`timescale 1ns/1ns
module testbench();
	wire[15:0] x, y, s;
	wire p, g, cin, cout;
	testAdder test(x, y, s, cin, cout);	
	add16 pfa1 (cout, s, p, g, x, y, cin);
endmodule

module testAdder(a, b, s, cin, cout);
	input [15:0] s, p, g;
	input cout;
	output [15:0] a, b;
	output cin;
	reg [15:0] a, b;
	reg cin;
	initial begin
		$monitor($time,,"a = %d, b = %d, cin = %b, s = %d, cout = %b", a, b, cin, s, cout);
	#10 a = 16687; b = 3597; cin = 1;
#10 a = 14642; b = 25400; cin = 1;
#10 a = 29923; b = 60414; cin = 1;
#10 a = 18974; b = 64900; cin = 1;
#10 a = 3642; b = 67258; cin = 0;
#10 a = 34114; b = 54843; cin = 0;
#10 a = 15634; b = 49945; cin = 1;
#10 a = 33270; b = 19719; cin = 1;
#10 a = 32910; b = 60722; cin = 0;
#10 a = 10070; b = 50511; cin = 1;
#10 a = 5154; b = 67198; cin = 1;
#10 a = 31951; b = 58193; cin = 1;
#10 a = 8309; b = 18116; cin = 1;
#10 a = 38534; b = 37091; cin = 1;
#10 a = 25539; b = 17085; cin = 0;
#10 a = 33313; b = 27551; cin = 1;
#10 a = 44077; b = 43186; cin = 0;
#10 a = 40436; b = 6456; cin = 1;
#10 a = 9757; b = 15719; cin = 1;
#10 a = 10837; b = 25789; cin = 1;
#10 a = 58799; b = 7296; cin = 1;
#10 a = 40358; b = 15599; cin = 0;
#10 a = 47317; b = 260; cin = 1;
#10 a = 67394; b = 38794; cin = 0;
#10 a = 36019; b = 64333; cin = 1;
#10 a = 48255; b = 27646; cin = 1;
#10 a = 21686; b = 48075; cin = 1;
#10 a = 45062; b = 64863; cin = 1;
#10 a = 64509; b = 4621; cin = 0;
#10 a = 4679; b = 61810; cin = 0;
#10 a = 19008; b = 26961; cin = 0;
#10 a = 53239; b = 67319; cin = 1;
#10 a = 5664; b = 20988; cin = 0;
#10 a = 22557; b = 18382; cin = 0;
#10 a = 6541; b = 54402; cin = 0;
#10 a = 53962; b = 9009; cin = 0;
#10 a = 58935; b = 7048; cin = 0;
#10 a = 37094; b = 28462; cin = 1;
#10 a = 68062; b = 22972; cin = 0;
#10 a = 21100; b = 27651; cin = 1;
#10 a = 46280; b = 23011; cin = 0;
#10 a = 8756; b = 52602; cin = 0;
#10 a = 33184; b = 58266; cin = 0;
#10 a = 57872; b = 10823; cin = 1;
#10 a = 51354; b = 63716; cin = 1;
#10 a = 39170; b = 47679; cin = 0;
#10 a = 7337; b = 36614; cin = 0;
#10 a = 47227; b = 50061; cin = 1;
#10 a = 58332; b = 24475; cin = 1;
#10 a = 50411; b = 21927; cin = 0;
#10 a = 10652; b = 68208; cin = 1;
#10 a = 67854; b = 6964; cin = 1;
#10 a = 52376; b = 16500; cin = 0;
#10 a = 34239; b = 4372; cin = 1;
#10 a = 34484; b = 55727; cin = 0;
#10 a = 65483; b = 1249; cin = 1;
#10 a = 35491; b = 8586; cin = 1;
#10 a = 35252; b = 55813; cin = 0;
#10 a = 63475; b = 20498; cin = 1;
#10 a = 21022; b = 909; cin = 1;
#10 a = 6220; b = 11561; cin = 1;
#10 a = 60781; b = 9415; cin = 1;
#10 a = 27944; b = 38144; cin = 0;
#10 a = 29726; b = 2383; cin = 0;
#10 a = 18684; b = 36867; cin = 1;
#10 a = 47710; b = 32350; cin = 1;
#10 a = 54415; b = 44193; cin = 1;
#10 a = 4086; b = 9445; cin = 1;
#10 a = 3819; b = 49272; cin = 1;
#10 a = 4378; b = 294; cin = 0;
#10 a = 26865; b = 6514; cin = 1;
#10 a = 47560; b = 43647; cin = 0;
#10 a = 51572; b = 47944; cin = 0;
#10 a = 48436; b = 7670; cin = 1;
#10 a = 49672; b = 2706; cin = 0;
#10 a = 36636; b = 26768; cin = 0;
#10 a = 1201; b = 11183; cin = 0;
#10 a = 68000; b = 15270; cin = 1;
#10 a = 3317; b = 65441; cin = 0;
#10 a = 29132; b = 69819; cin = 0;
#10 a = 32208; b = 3037; cin = 1;
#10 a = 23197; b = 50597; cin = 0;
#10 a = 23602; b = 8521; cin = 0;
#10 a = 38502; b = 33309; cin = 1;
#10 a = 32138; b = 12982; cin = 1;
#10 a = 62640; b = 25970; cin = 0;
#10 a = 55493; b = 27171; cin = 1;
#10 a = 68891; b = 1523; cin = 1;
#10 a = 68086; b = 4841; cin = 0;
#10 a = 46554; b = 10325; cin = 0;
#10 a = 25317; b = 42534; cin = 1;
#10 a = 56946; b = 65731; cin = 0;
#10 a = 62222; b = 65685; cin = 0;
#10 a = 45443; b = 10540; cin = 1;
#10 a = 59038; b = 42678; cin = 1;
#10 a = 28987; b = 11670; cin = 1;
#10 a = 2057; b = 43515; cin = 0;
#10 a = 32663; b = 42406; cin = 0;
#10 a = 8538; b = 16845; cin = 1;
#10 a = 49855; b = 63399; cin = 0;
#10 a = 67343; b = 18716; cin = 0;
#10 a = 17868; b = 52014; cin = 0;
#10 a = 65342; b = 20589; cin = 1;
#10 a = 27690; b = 42384; cin = 1;
#10 a = 23348; b = 31422; cin = 1;
#10 a = 31987; b = 36761; cin = 0;
#10 a = 42949; b = 38819; cin = 1;
#10 a = 11081; b = 47834; cin = 0;
#10 a = 27089; b = 56372; cin = 1;
#10 a = 47938; b = 36227; cin = 0;
#10 a = 9113; b = 9922; cin = 1;
#10 a = 12821; b = 4142; cin = 1;
#10 a = 58613; b = 45837; cin = 0;
#10 a = 6443; b = 3527; cin = 0;
#10 a = 34812; b = 3227; cin = 0;
#10 a = 12212; b = 11567; cin = 0;
#10 a = 24930; b = 54516; cin = 1;
#10 a = 57515; b = 41949; cin = 1;
#10 a = 38859; b = 69039; cin = 1;
#10 a = 37048; b = 46977; cin = 1;
#10 a = 28637; b = 32442; cin = 1;
#10 a = 15294; b = 45264; cin = 0;
#10 a = 53965; b = 10229; cin = 1;
#10 a = 43226; b = 63024; cin = 0;
#10 a = 51222; b = 27837; cin = 0;
#10 a = 44289; b = 40049; cin = 1;
#10 a = 4117; b = 41331; cin = 1;
#10 a = 25468; b = 5198; cin = 0;
#10 a = 48301; b = 20410; cin = 1;
#10 a = 33858; b = 57458; cin = 1;
#10 a = 55643; b = 62447; cin = 1;
#10 a = 40055; b = 7741; cin = 1;
#10 a = 52257; b = 38059; cin = 1;
#10 a = 16648; b = 11285; cin = 1;
#10 a = 30918; b = 62507; cin = 0;
#10 a = 2064; b = 13148; cin = 1;
#10 a = 31129; b = 63617; cin = 0;
#10 a = 21062; b = 19085; cin = 1;
#10 a = 52945; b = 67386; cin = 1;
#10 a = 60218; b = 7597; cin = 1;
#10 a = 20821; b = 39592; cin = 1;
#10 a = 13867; b = 9647; cin = 0;
#10 a = 28528; b = 38256; cin = 1;
#10 a = 29771; b = 54904; cin = 0;
#10 a = 24039; b = 15823; cin = 0;
#10 a = 22495; b = 64239; cin = 0;
#10 a = 37353; b = 25369; cin = 0;
#10 a = 69893; b = 22783; cin = 1;
#10 a = 37632; b = 5728; cin = 0;
#10 a = 2133; b = 65947; cin = 1;
#10 a = 445; b = 16768; cin = 1;
#10 a = 61204; b = 6987; cin = 1;
#10 a = 59704; b = 35516; cin = 1;
#10 a = 2616; b = 65287; cin = 0;
#10 a = 26812; b = 65678; cin = 1;
#10 a = 19868; b = 64526; cin = 0;
#10 a = 26073; b = 8231; cin = 1;
#10 a = 25895; b = 8124; cin = 1;
#10 a = 21154; b = 22109; cin = 1;
#10 a = 13800; b = 594; cin = 0;
#10 a = 60395; b = 47391; cin = 1;
#10 a = 6583; b = 38595; cin = 0;
#10 a = 32418; b = 4652; cin = 0;
#10 a = 26509; b = 7268; cin = 0;
#10 a = 51857; b = 10432; cin = 0;
#10 a = 23028; b = 30301; cin = 0;
#10 a = 34791; b = 32726; cin = 1;
#10 a = 1922; b = 34973; cin = 0;
#10 a = 38189; b = 56127; cin = 1;
#10 a = 10185; b = 46280; cin = 1;
#10 a = 24479; b = 13027; cin = 1;
#10 a = 31894; b = 19610; cin = 0;
#10 a = 46297; b = 28380; cin = 0;
#10 a = 2567; b = 54890; cin = 0;
#10 a = 24125; b = 36747; cin = 1;
#10 a = 17714; b = 36128; cin = 0;
#10 a = 5828; b = 919; cin = 0;
#10 a = 48526; b = 49193; cin = 1;
#10 a = 29348; b = 63735; cin = 0;
#10 a = 8631; b = 3920; cin = 0;
#10 a = 58508; b = 4751; cin = 0;
#10 a = 62129; b = 36646; cin = 0;
#10 a = 34346; b = 59295; cin = 1;
#10 a = 11214; b = 61862; cin = 1;
#10 a = 41703; b = 62340; cin = 0;
#10 a = 58976; b = 10054; cin = 0;
#10 a = 36550; b = 62234; cin = 1;
#10 a = 23202; b = 40760; cin = 1;
#10 a = 44827; b = 46460; cin = 0;
#10 a = 28931; b = 55091; cin = 0;
#10 a = 35668; b = 19952; cin = 1;
#10 a = 31784; b = 12081; cin = 1;
#10 a = 47510; b = 46427; cin = 0;
#10 a = 21617; b = 57642; cin = 1;
#10 a = 3318; b = 5697; cin = 1;
#10 a = 21767; b = 64673; cin = 1;
#10 a = 52695; b = 7575; cin = 1;
#10 a = 14543; b = 30777; cin = 0;
#10 a = 1936; b = 5604; cin = 0;
#10 a = 53064; b = 34535; cin = 0;
#10 a = 14464; b = 46555; cin = 0;
#10 a = 50615; b = 8339; cin = 1;
#10 a = 6117; b = 55850; cin = 1;
#10 a = 20913; b = 53819; cin = 1;
#10 a = 27572; b = 33490; cin = 0;
#10 a = 2923; b = 55257; cin = 1;
#10 a = 58328; b = 37952; cin = 0;
#10 a = 12320; b = 28847; cin = 1;
#10 a = 7072; b = 30783; cin = 1;
#10 a = 24636; b = 60199; cin = 0;
#10 a = 50940; b = 51015; cin = 0;
#10 a = 3548; b = 31631; cin = 1;
#10 a = 38238; b = 14100; cin = 1;
#10 a = 49355; b = 35013; cin = 1;
#10 a = 24466; b = 38938; cin = 1;
#10 a = 5274; b = 41861; cin = 0;
#10 a = 27107; b = 6542; cin = 0;
#10 a = 56515; b = 65214; cin = 0;
#10 a = 46700; b = 48638; cin = 1;
#10 a = 18841; b = 3274; cin = 1;
#10 a = 1869; b = 30567; cin = 0;
#10 a = 31453; b = 34115; cin = 1;
#10 a = 69377; b = 48705; cin = 1;
#10 a = 45854; b = 28060; cin = 1;
#10 a = 6151; b = 52526; cin = 1;
#10 a = 69938; b = 34152; cin = 0;
#10 a = 1686; b = 37611; cin = 0;
#10 a = 41387; b = 478; cin = 0;
#10 a = 39935; b = 23530; cin = 0;
#10 a = 21970; b = 42371; cin = 1;
#10 a = 64205; b = 44241; cin = 0;
#10 a = 17456; b = 5694; cin = 1;
#10 a = 48689; b = 51423; cin = 1;
#10 a = 24023; b = 27278; cin = 1;
#10 a = 10722; b = 9781; cin = 0;
#10 a = 36359; b = 56072; cin = 0;
#10 a = 10209; b = 57758; cin = 0;
#10 a = 36954; b = 29145; cin = 0;
#10 a = 58912; b = 45432; cin = 1;
#10 a = 59509; b = 67403; cin = 0;
#10 a = 63380; b = 61608; cin = 1;
#10 a = 27818; b = 9064; cin = 0;
#10 a = 2723; b = 57754; cin = 1;
#10 a = 26334; b = 58129; cin = 1;
#10 a = 54358; b = 68851; cin = 1;
#10 a = 41260; b = 11562; cin = 1;
#10 a = 62314; b = 21771; cin = 1;
#10 a = 50980; b = 58725; cin = 1;
#10 a = 16477; b = 23990; cin = 1;
#10 a = 5504; b = 13499; cin = 0;
#10 a = 13254; b = 53231; cin = 1;
#10 a = 65246; b = 57401; cin = 1;
#10 a = 5636; b = 60124; cin = 1;
#10 a = 67449; b = 62811; cin = 0;
#10 a = 62893; b = 23521; cin = 1;
#10 a = 21766; b = 64781; cin = 1;
#10 a = 13063; b = 57095; cin = 1;
#10 a = 62118; b = 14428; cin = 0;
#10 a = 46671; b = 7257; cin = 0;
#10 a = 6657; b = 59113; cin = 1;
#10 a = 34045; b = 2367; cin = 0;
#10 a = 53042; b = 43965; cin = 1;
#10 a = 57456; b = 49601; cin = 0;
#10 a = 49623; b = 23403; cin = 1;
#10 a = 6272; b = 16296; cin = 0;
#10 a = 8123; b = 14414; cin = 1;
#10 a = 21537; b = 3829; cin = 0;
#10 a = 56722; b = 42299; cin = 0;
#10 a = 56984; b = 18971; cin = 1;
#10 a = 57589; b = 25628; cin = 0;
#10 a = 1692; b = 59673; cin = 0;
#10 a = 69027; b = 19068; cin = 1;
#10 a = 53762; b = 6524; cin = 1;
#10 a = 4974; b = 32499; cin = 0;
#10 a = 65349; b = 15123; cin = 0;
#10 a = 9245; b = 23247; cin = 0;
#10 a = 64274; b = 44784; cin = 1;
#10 a = 12751; b = 7858; cin = 0;
#10 a = 22007; b = 64842; cin = 1;
#10 a = 38521; b = 52431; cin = 1;
#10 a = 44147; b = 54124; cin = 1;
#10 a = 28493; b = 29503; cin = 1;
#10 a = 56805; b = 13265; cin = 1;
#10 a = 41070; b = 18240; cin = 0;
#10 a = 48738; b = 13589; cin = 0;
#10 a = 2702; b = 69187; cin = 1;
#10 a = 17432; b = 63461; cin = 1;
#10 a = 35991; b = 52564; cin = 1;
#10 a = 3201; b = 4572; cin = 1;
#10 a = 59383; b = 19445; cin = 1;
#10 a = 47544; b = 63592; cin = 1;
#10 a = 1731; b = 68438; cin = 0;
#10 a = 44986; b = 55243; cin = 1;
#10 a = 24765; b = 26313; cin = 1;
#10 a = 13396; b = 51403; cin = 1;
#10 a = 17150; b = 54105; cin = 0;
#10 a = 44151; b = 47889; cin = 1;
#10 a = 22288; b = 60232; cin = 0;
#10 a = 8283; b = 63433; cin = 0;
#10 a = 35472; b = 29168; cin = 1;
#10 a = 45093; b = 6713; cin = 1;
#10 a = 61542; b = 8444; cin = 1;
#10 a = 61142; b = 53431; cin = 0;
#10 a = 4008; b = 54548; cin = 1;
#10 a = 57817; b = 44296; cin = 0;
#10 a = 55216; b = 61446; cin = 1;
#10 a = 28154; b = 11949; cin = 0;
#10 a = 64554; b = 34237; cin = 0;
#10 a = 59870; b = 18872; cin = 0;
#10 a = 36110; b = 54345; cin = 0;
#10 a = 31795; b = 5790; cin = 1;
#10 a = 21072; b = 67333; cin = 0;
#10 a = 8788; b = 34827; cin = 1;
#10 a = 28098; b = 15187; cin = 1;
#10 a = 50074; b = 3005; cin = 0;
#10 a = 7100; b = 58221; cin = 0;
#10 a = 40936; b = 16376; cin = 0;
#10 a = 52660; b = 57282; cin = 1;
#10 a = 30969; b = 23504; cin = 0;
#10 a = 2711; b = 59614; cin = 1;
#10 a = 3621; b = 21409; cin = 1;
#10 a = 33949; b = 42481; cin = 0;
#10 a = 26369; b = 27621; cin = 0;
#10 a = 24924; b = 32072; cin = 1;
#10 a = 8027; b = 12146; cin = 0;
#10 a = 11779; b = 65598; cin = 0;
#10 a = 30626; b = 12886; cin = 0;
#10 a = 37774; b = 65547; cin = 0;
#10 a = 55511; b = 26516; cin = 0;
#10 a = 22121; b = 29227; cin = 0;
#10 a = 43076; b = 9200; cin = 1;
#10 a = 22526; b = 43149; cin = 0;
#10 a = 69308; b = 45870; cin = 0;
#10 a = 10918; b = 47146; cin = 0;
#10 a = 37716; b = 55174; cin = 0;
#10 a = 43870; b = 66953; cin = 0;
#10 a = 38246; b = 3931; cin = 1;
#10 a = 25350; b = 18057; cin = 0;
#10 a = 46088; b = 49921; cin = 0;
#10 a = 20330; b = 2042; cin = 1;
#10 a = 54186; b = 21471; cin = 1;
#10 a = 39451; b = 43997; cin = 1;
#10 a = 19902; b = 43305; cin = 1;
#10 a = 27974; b = 54224; cin = 0;
#10 a = 44470; b = 68292; cin = 0;
#10 a = 3112; b = 42162; cin = 1;
#10 a = 50056; b = 56761; cin = 1;
#10 a = 63535; b = 12111; cin = 0;
#10 a = 48913; b = 34552; cin = 1;
#10 a = 37159; b = 54882; cin = 0;
#10 a = 54632; b = 39069; cin = 1;
#10 a = 34010; b = 54872; cin = 0;
#10 a = 56537; b = 51126; cin = 1;
#10 a = 7638; b = 9100; cin = 1;
#10 a = 29534; b = 29922; cin = 1;
#10 a = 12956; b = 9386; cin = 0;
#10 a = 39684; b = 59443; cin = 1;
#10 a = 46695; b = 29330; cin = 0;
#10 a = 1763; b = 54596; cin = 0;
#10 a = 53105; b = 21755; cin = 1;
#10 a = 60137; b = 52740; cin = 0;
#10 a = 64992; b = 16750; cin = 0;
#10 a = 20196; b = 49639; cin = 1;
#10 a = 18705; b = 57277; cin = 1;
#10 a = 1439; b = 63164; cin = 0;
#10 a = 28816; b = 6120; cin = 0;
#10 a = 28356; b = 45804; cin = 1;
#10 a = 14657; b = 22499; cin = 0;
#10 a = 59422; b = 615; cin = 0;
#10 a = 68738; b = 53720; cin = 1;
#10 a = 39289; b = 20209; cin = 1;
#10 a = 1613; b = 61553; cin = 1;
#10 a = 18810; b = 11749; cin = 0;
#10 a = 17133; b = 30454; cin = 0;
#10 a = 908; b = 8245; cin = 0;
#10 a = 14606; b = 37062; cin = 0;
#10 a = 37691; b = 65418; cin = 1;
#10 a = 26570; b = 10076; cin = 0;
#10 a = 44780; b = 69498; cin = 1;
#10 a = 47586; b = 44588; cin = 1;
#10 a = 48500; b = 60230; cin = 0;
#10 a = 8505; b = 61843; cin = 1;
#10 a = 55261; b = 10653; cin = 0;
#10 a = 34359; b = 27786; cin = 1;
#10 a = 735; b = 28695; cin = 0;
#10 a = 30275; b = 19653; cin = 0;
#10 a = 42288; b = 33696; cin = 1;
#10 a = 6457; b = 60267; cin = 1;
#10 a = 63125; b = 11399; cin = 1;
#10 a = 26761; b = 35338; cin = 1;
#10 a = 20468; b = 13838; cin = 1;
#10 a = 58033; b = 68695; cin = 1;
#10 a = 63502; b = 53956; cin = 0;
#10 a = 10721; b = 18316; cin = 1;
#10 a = 34746; b = 19051; cin = 0;
#10 a = 67016; b = 25679; cin = 1;
#10 a = 66349; b = 67967; cin = 0;
#10 a = 61100; b = 50776; cin = 1;
#10 a = 42279; b = 43901; cin = 0;
#10 a = 22956; b = 47014; cin = 0;
#10 a = 48221; b = 67483; cin = 0;
#10 a = 63717; b = 31868; cin = 0;
#10 a = 1056; b = 1722; cin = 0;
#10 a = 65400; b = 12443; cin = 0;
#10 a = 17531; b = 23541; cin = 0;
#10 a = 44709; b = 66910; cin = 1;
#10 a = 21541; b = 63259; cin = 0;
#10 a = 32069; b = 30711; cin = 0;
#10 a = 55568; b = 2990; cin = 1;
#10 a = 44114; b = 25946; cin = 0;
#10 a = 67999; b = 50519; cin = 1;
#10 a = 12073; b = 44236; cin = 1;
#10 a = 1195; b = 21644; cin = 1;
#10 a = 44274; b = 17045; cin = 1;
#10 a = 35668; b = 34576; cin = 0;
#10 a = 68818; b = 9286; cin = 0;
#10 a = 57647; b = 30827; cin = 1;
#10 a = 20795; b = 39248; cin = 0;
#10 a = 11071; b = 24816; cin = 0;
#10 a = 45249; b = 45282; cin = 0;
#10 a = 32793; b = 19633; cin = 0;
#10 a = 64172; b = 8059; cin = 0;
#10 a = 33771; b = 9254; cin = 1;
#10 a = 28740; b = 53528; cin = 0;
#10 a = 58857; b = 19197; cin = 0;
#10 a = 42516; b = 64367; cin = 0;
#10 a = 69436; b = 28367; cin = 1;
#10 a = 19616; b = 25514; cin = 1;
#10 a = 506; b = 36586; cin = 1;
#10 a = 7091; b = 58187; cin = 0;
#10 a = 39621; b = 20980; cin = 1;
#10 a = 52671; b = 61504; cin = 0;
#10 a = 39958; b = 25275; cin = 1;
#10 a = 25241; b = 30367; cin = 1;
#10 a = 3921; b = 65577; cin = 0;
#10 a = 40825; b = 14445; cin = 0;
#10 a = 39720; b = 13881; cin = 1;
#10 a = 69441; b = 33497; cin = 1;
#10 a = 44763; b = 10356; cin = 1;
#10 a = 67604; b = 17447; cin = 0;
#10 a = 19376; b = 57068; cin = 0;
#10 a = 37134; b = 39740; cin = 0;
#10 a = 62950; b = 56050; cin = 1;
#10 a = 28021; b = 57643; cin = 1;
#10 a = 46621; b = 61564; cin = 0;
#10 a = 14417; b = 8741; cin = 1;
#10 a = 69285; b = 48461; cin = 0;
#10 a = 36168; b = 24255; cin = 0;
#10 a = 28566; b = 45370; cin = 0;
#10 a = 33901; b = 42974; cin = 1;
#10 a = 27424; b = 38703; cin = 1;
#10 a = 41926; b = 5837; cin = 1;
#10 a = 637; b = 45139; cin = 1;
#10 a = 54622; b = 3161; cin = 0;
#10 a = 68975; b = 49782; cin = 0;
#10 a = 31609; b = 40551; cin = 0;
#10 a = 32336; b = 39837; cin = 1;
#10 a = 23297; b = 6005; cin = 0;
#10 a = 47755; b = 10923; cin = 0;
#10 a = 58921; b = 21177; cin = 1;
#10 a = 17534; b = 48601; cin = 0;
#10 a = 9567; b = 66879; cin = 1;
#10 a = 41341; b = 67516; cin = 0;
#10 a = 35516; b = 52139; cin = 1;
#10 a = 63687; b = 27466; cin = 1;
#10 a = 13421; b = 35428; cin = 1;
#10 a = 18249; b = 67764; cin = 0;
#10 a = 47891; b = 67413; cin = 1;
#10 a = 31787; b = 45168; cin = 1;
#10 a = 37406; b = 10441; cin = 0;
#10 a = 15999; b = 27975; cin = 1;
#10 a = 33295; b = 37543; cin = 0;
#10 a = 32780; b = 55236; cin = 1;
#10 a = 7404; b = 67104; cin = 0;
#10 a = 55190; b = 60791; cin = 0;
#10 a = 12757; b = 50565; cin = 0;
#10 a = 57228; b = 45166; cin = 1;
#10 a = 1536; b = 69409; cin = 0;
#10 a = 68202; b = 7549; cin = 1;
#10 a = 52143; b = 44955; cin = 0;
#10 a = 57261; b = 37306; cin = 0;
#10 a = 40980; b = 601; cin = 1;
#10 a = 67930; b = 33381; cin = 1;
#10 a = 45101; b = 40785; cin = 1;
#10 a = 4411; b = 2327; cin = 1;
#10 a = 37540; b = 15085; cin = 0;
#10 a = 36096; b = 48665; cin = 0;
#10 a = 8769; b = 50202; cin = 0;
#10 a = 48856; b = 48404; cin = 1;
#10 a = 40463; b = 30547; cin = 0;
#10 a = 18863; b = 64160; cin = 0;
#10 a = 25239; b = 35140; cin = 1;
#10 a = 69158; b = 9422; cin = 0;
#10 a = 4665; b = 54524; cin = 1;
#10 a = 7277; b = 35287; cin = 1;
#10 a = 47032; b = 2827; cin = 0;
#10 a = 67352; b = 38924; cin = 1;
#10 a = 62838; b = 24045; cin = 1;
#10 a = 34086; b = 2901; cin = 1;
#10 a = 36531; b = 19716; cin = 0;
#10 a = 36635; b = 38580; cin = 0;
#10 a = 27693; b = 63819; cin = 0;
#10 a = 65704; b = 39330; cin = 1;
#10 a = 43448; b = 20347; cin = 1;
#10 a = 38330; b = 27624; cin = 0;
#10 a = 35539; b = 4656; cin = 0;
#10 a = 47833; b = 2008; cin = 0;
#10 a = 15144; b = 41199; cin = 1;
#10 a = 32658; b = 5285; cin = 1;
#10 a = 4927; b = 18169; cin = 1;
#10 a = 54096; b = 54804; cin = 1;
#10 a = 3776; b = 12498; cin = 1;
#10 a = 12245; b = 54554; cin = 1;
#10 a = 52840; b = 28003; cin = 0;
#10 a = 7959; b = 66333; cin = 1;
#10 a = 68365; b = 8224; cin = 1;
#10 a = 37951; b = 56057; cin = 0;
#10 a = 46461; b = 47553; cin = 1;
#10 a = 9017; b = 56563; cin = 0;
#10 a = 20826; b = 61491; cin = 1;
#10 a = 28703; b = 21939; cin = 0;
#10 a = 28809; b = 25715; cin = 0;
#10 a = 45438; b = 14312; cin = 0;
#10 a = 31397; b = 43504; cin = 1;
#10 a = 37703; b = 51463; cin = 0;
#10 a = 1634; b = 26181; cin = 0;
#10 a = 62926; b = 40484; cin = 1;
#10 a = 56226; b = 16946; cin = 1;
#10 a = 20725; b = 2315; cin = 0;
#10 a = 36861; b = 69493; cin = 1;
#10 a = 47519; b = 28196; cin = 0;
#10 a = 66629; b = 33357; cin = 0;
#10 a = 50941; b = 8795; cin = 0;
#10 a = 19807; b = 40192; cin = 1;
#10 a = 16677; b = 7896; cin = 0;
#10 a = 32583; b = 55882; cin = 1;
#10 a = 56714; b = 48808; cin = 0;
#10 a = 43253; b = 11386; cin = 0;
#10 a = 7346; b = 8463; cin = 1;
#10 a = 28003; b = 45325; cin = 0;
#10 a = 16502; b = 22844; cin = 0;
#10 a = 3293; b = 65825; cin = 0;
#10 a = 62151; b = 46766; cin = 1;
#10 a = 41673; b = 66573; cin = 0;
#10 a = 64700; b = 59602; cin = 0;
#10 a = 45543; b = 22186; cin = 0;
#10 a = 52566; b = 55252; cin = 1;
#10 a = 30074; b = 28505; cin = 1;
#10 a = 880; b = 35852; cin = 1;
#10 a = 20353; b = 40207; cin = 0;
#10 a = 15671; b = 33061; cin = 0;
#10 a = 39186; b = 12706; cin = 1;
#10 a = 26058; b = 51209; cin = 1;
#10 a = 68077; b = 69235; cin = 0;
#10 a = 56641; b = 63935; cin = 1;
#10 a = 29453; b = 39478; cin = 1;
#10 a = 58148; b = 22045; cin = 1;
#10 a = 18355; b = 28471; cin = 0;
#10 a = 13596; b = 5704; cin = 0;
#10 a = 63653; b = 2409; cin = 1;
#10 a = 65387; b = 18081; cin = 1;
#10 a = 19965; b = 57267; cin = 1;
#10 a = 16720; b = 13325; cin = 1;
#10 a = 36593; b = 57754; cin = 0;
#10 a = 29392; b = 20748; cin = 1;
#10 a = 35441; b = 50201; cin = 0;
#10 a = 16380; b = 14701; cin = 1;
#10 a = 52571; b = 33056; cin = 0;
#10 a = 23619; b = 23005; cin = 0;
#10 a = 30520; b = 63010; cin = 0;
#10 a = 30331; b = 58398; cin = 1;
#10 a = 16852; b = 54715; cin = 0;
#10 a = 62432; b = 47788; cin = 1;
#10 a = 19221; b = 60733; cin = 1;
#10 a = 21597; b = 20125; cin = 1;
#10 a = 17908; b = 55566; cin = 1;
#10 a = 53698; b = 48298; cin = 0;
#10 a = 17885; b = 30869; cin = 1;
#10 a = 56896; b = 30841; cin = 0;
#10 a = 31610; b = 37713; cin = 0;
#10 a = 55086; b = 68044; cin = 0;
#10 a = 50291; b = 14897; cin = 0;
#10 a = 9115; b = 53681; cin = 0;
#10 a = 27616; b = 49254; cin = 1;
#10 a = 33872; b = 851; cin = 1;
#10 a = 60875; b = 18759; cin = 1;
#10 a = 44432; b = 2458; cin = 0;
#10 a = 42691; b = 66695; cin = 1;
#10 a = 50358; b = 29943; cin = 0;
#10 a = 57382; b = 37906; cin = 1;
#10 a = 57416; b = 22992; cin = 0;
#10 a = 22201; b = 3284; cin = 1;
#10 a = 41701; b = 58751; cin = 0;
#10 a = 38989; b = 16368; cin = 0;
#10 a = 3362; b = 50240; cin = 1;
#10 a = 57861; b = 17467; cin = 0;
#10 a = 27927; b = 61900; cin = 0;
#10 a = 22643; b = 10943; cin = 0;
#10 a = 24580; b = 61301; cin = 1;
#10 a = 57359; b = 48683; cin = 1;
#10 a = 57850; b = 12451; cin = 0;
#10 a = 56386; b = 34652; cin = 0;
#10 a = 46171; b = 6353; cin = 1;
#10 a = 19637; b = 45342; cin = 1;
#10 a = 42357; b = 25057; cin = 1;
#10 a = 65928; b = 12918; cin = 1;
#10 a = 38259; b = 40845; cin = 1;
#10 a = 35751; b = 39840; cin = 0;
#10 a = 29939; b = 64421; cin = 1;
#10 a = 30423; b = 51780; cin = 0;
#10 a = 68812; b = 39630; cin = 1;
#10 a = 36546; b = 2369; cin = 0;
#10 a = 53916; b = 48540; cin = 1;
#10 a = 60038; b = 68178; cin = 0;
#10 a = 58879; b = 40535; cin = 1;
#10 a = 37961; b = 12816; cin = 1;
#10 a = 34510; b = 51075; cin = 1;
#10 a = 69311; b = 63178; cin = 1;
#10 a = 45055; b = 23118; cin = 0;
#10 a = 12100; b = 29893; cin = 0;
#10 a = 50532; b = 5057; cin = 1;
#10 a = 55063; b = 41604; cin = 0;
#10 a = 599; b = 1872; cin = 0;
#10 a = 46137; b = 61910; cin = 0;
#10 a = 19721; b = 50790; cin = 0;
#10 a = 18362; b = 18751; cin = 0;
#10 a = 29921; b = 29613; cin = 1;
#10 a = 58678; b = 28924; cin = 1;
#10 a = 33628; b = 3979; cin = 1;
#10 a = 2998; b = 62431; cin = 0;
#10 a = 501; b = 19315; cin = 0;
#10 a = 37634; b = 4378; cin = 0;
#10 a = 53488; b = 4978; cin = 0;
#10 a = 47882; b = 27467; cin = 1;
#10 a = 40455; b = 23540; cin = 1;
#10 a = 49915; b = 41902; cin = 0;
#10 a = 2191; b = 48175; cin = 1;
#10 a = 51894; b = 13206; cin = 1;
#10 a = 24775; b = 46834; cin = 0;
#10 a = 43479; b = 26184; cin = 1;
#10 a = 45723; b = 26685; cin = 0;
#10 a = 29377; b = 64319; cin = 0;
#10 a = 54635; b = 24159; cin = 0;
#10 a = 11766; b = 2042; cin = 1;
#10 a = 7159; b = 42497; cin = 1;
#10 a = 29694; b = 22412; cin = 1;
#10 a = 47332; b = 955; cin = 1;
#10 a = 24583; b = 52849; cin = 1;
#10 a = 7110; b = 53976; cin = 1;
#10 a = 39968; b = 27455; cin = 1;
#10 a = 41609; b = 49531; cin = 1;
#10 a = 16213; b = 8908; cin = 0;
#10 a = 17899; b = 63544; cin = 0;
#10 a = 24564; b = 5310; cin = 0;
#10 a = 35047; b = 58821; cin = 1;
#10 a = 45423; b = 18515; cin = 1;
#10 a = 27700; b = 42199; cin = 0;
#10 a = 58153; b = 43134; cin = 1;
#10 a = 8164; b = 50244; cin = 1;
#10 a = 5009; b = 66564; cin = 1;
#10 a = 4391; b = 38173; cin = 0;
#10 a = 30458; b = 30738; cin = 0;
#10 a = 27196; b = 48637; cin = 0;
#10 a = 48094; b = 49553; cin = 0;
#10 a = 1034; b = 14601; cin = 1;
#10 a = 42823; b = 60024; cin = 0;
#10 a = 13376; b = 17724; cin = 1;
#10 a = 8532; b = 52230; cin = 1;
#10 a = 9241; b = 60394; cin = 1;
#10 a = 63927; b = 65404; cin = 1;
#10 a = 52420; b = 46147; cin = 0;
#10 a = 44092; b = 6605; cin = 0;
#10 a = 67376; b = 10153; cin = 0;
#10 a = 37853; b = 58248; cin = 1;
#10 a = 36343; b = 35634; cin = 0;
#10 a = 23655; b = 54810; cin = 0;
#10 a = 5833; b = 68186; cin = 1;
#10 a = 30211; b = 53071; cin = 1;
#10 a = 4074; b = 62312; cin = 1;
#10 a = 28182; b = 56239; cin = 1;
#10 a = 25205; b = 38659; cin = 0;
#10 a = 60402; b = 59103; cin = 1;
#10 a = 32688; b = 32832; cin = 1;
#10 a = 53612; b = 685; cin = 1;
#10 a = 54090; b = 13380; cin = 1;
#10 a = 45520; b = 37035; cin = 1;
#10 a = 3327; b = 19221; cin = 0;
#10 a = 25210; b = 25784; cin = 1;
#10 a = 5675; b = 29858; cin = 1;
#10 a = 182; b = 34392; cin = 1;
#10 a = 12798; b = 59598; cin = 0;
#10 a = 1560; b = 26352; cin = 0;
#10 a = 66928; b = 59040; cin = 0;
#10 a = 48801; b = 19005; cin = 1;
#10 a = 18922; b = 49447; cin = 1;
#10 a = 1029; b = 24967; cin = 1;
#10 a = 14299; b = 4646; cin = 0;
#10 a = 25755; b = 6208; cin = 0;
#10 a = 20282; b = 11883; cin = 0;
#10 a = 7121; b = 58418; cin = 1;
#10 a = 2904; b = 47568; cin = 1;
#10 a = 37347; b = 49128; cin = 1;
#10 a = 13597; b = 22408; cin = 1;
#10 a = 46327; b = 47561; cin = 0;
#10 a = 32446; b = 66483; cin = 1;
#10 a = 31945; b = 43865; cin = 1;
#10 a = 44832; b = 58164; cin = 1;
#10 a = 6940; b = 13919; cin = 0;
#10 a = 64832; b = 10553; cin = 1;
#10 a = 12583; b = 17674; cin = 1;
#10 a = 41078; b = 66931; cin = 1;
#10 a = 59171; b = 10630; cin = 0;
#10 a = 9968; b = 24227; cin = 0;
#10 a = 66157; b = 46906; cin = 0;
#10 a = 1352; b = 9352; cin = 1;
#10 a = 32345; b = 17649; cin = 0;
#10 a = 18306; b = 62482; cin = 0;
#10 a = 55266; b = 69422; cin = 1;
#10 a = 4786; b = 64255; cin = 0;
#10 a = 36189; b = 53190; cin = 1;
#10 a = 8715; b = 24268; cin = 0;
#10 a = 28808; b = 59791; cin = 0;
#10 a = 4382; b = 69759; cin = 1;
#10 a = 48717; b = 42268; cin = 1;
#10 a = 613; b = 43620; cin = 1;
#10 a = 18992; b = 5966; cin = 0;
#10 a = 33941; b = 624; cin = 0;
#10 a = 60701; b = 55890; cin = 1;
#10 a = 54085; b = 60676; cin = 0;
#10 a = 58021; b = 3218; cin = 0;
#10 a = 55984; b = 11933; cin = 0;
#10 a = 50878; b = 17093; cin = 1;
#10 a = 56402; b = 67828; cin = 0;
#10 a = 16153; b = 46545; cin = 0;
#10 a = 69162; b = 47158; cin = 1;
#10 a = 61523; b = 42502; cin = 1;
#10 a = 47886; b = 6443; cin = 1;
#10 a = 26730; b = 43497; cin = 0;
#10 a = 4997; b = 3934; cin = 0;
#10 a = 223; b = 38307; cin = 0;
#10 a = 48639; b = 24292; cin = 1;
#10 a = 51323; b = 5170; cin = 1;
#10 a = 20150; b = 37925; cin = 1;
#10 a = 35088; b = 30430; cin = 0;
#10 a = 22295; b = 29593; cin = 0;
#10 a = 29474; b = 67468; cin = 0;
#10 a = 18971; b = 45354; cin = 0;
#10 a = 32740; b = 48437; cin = 1;
#10 a = 55104; b = 53434; cin = 1;
#10 a = 68145; b = 53658; cin = 0;
#10 a = 14403; b = 32297; cin = 0;
#10 a = 18947; b = 59973; cin = 1;
#10 a = 16936; b = 56475; cin = 0;
#10 a = 36401; b = 67916; cin = 0;
#10 a = 8763; b = 20211; cin = 1;
#10 a = 4635; b = 49685; cin = 0;
#10 a = 19361; b = 68656; cin = 0;
#10 a = 16883; b = 7748; cin = 1;
#10 a = 34254; b = 39205; cin = 0;
#10 a = 55559; b = 37350; cin = 0;
#10 a = 21524; b = 28105; cin = 1;
#10 a = 11780; b = 23404; cin = 0;
#10 a = 53559; b = 40340; cin = 0;
#10 a = 63263; b = 53093; cin = 0;
#10 a = 33398; b = 61856; cin = 1;
#10 a = 55829; b = 42843; cin = 0;
#10 a = 5729; b = 38557; cin = 0;
#10 a = 47336; b = 31792; cin = 0;
#10 a = 67379; b = 66047; cin = 1;
#10 a = 857; b = 27958; cin = 1;
#10 a = 10697; b = 49482; cin = 1;
#10 a = 52835; b = 61263; cin = 1;
#10 a = 61297; b = 44822; cin = 0;
#10 a = 32587; b = 14438; cin = 1;
#10 a = 25441; b = 47836; cin = 0;
#10 a = 14858; b = 10017; cin = 1;
#10 a = 30312; b = 15747; cin = 0;
#10 a = 20774; b = 63083; cin = 1;
#10 a = 65337; b = 60462; cin = 0;
#10 a = 9104; b = 37672; cin = 0;
#10 a = 60222; b = 48369; cin = 1;
#10 a = 22149; b = 7556; cin = 0;
#10 a = 31128; b = 45206; cin = 0;
#10 a = 56800; b = 7793; cin = 0;
#10 a = 65566; b = 9587; cin = 0;
#10 a = 42540; b = 797; cin = 0;
#10 a = 62357; b = 31110; cin = 1;
#10 a = 27084; b = 28236; cin = 0;
#10 a = 23603; b = 23573; cin = 0;
#10 a = 62521; b = 32678; cin = 0;
#10 a = 59397; b = 69252; cin = 0;
#10 a = 12108; b = 21401; cin = 0;
#10 a = 26082; b = 28881; cin = 0;
#10 a = 37583; b = 15682; cin = 0;
#10 a = 63521; b = 57600; cin = 1;
#10 a = 43648; b = 30140; cin = 0;
#10 a = 33792; b = 68849; cin = 0;
#10 a = 39683; b = 25933; cin = 1;
#10 a = 38657; b = 25888; cin = 0;
#10 a = 50797; b = 18409; cin = 0;
#10 a = 54258; b = 54159; cin = 0;
#10 a = 58792; b = 66267; cin = 1;
#10 a = 47234; b = 22350; cin = 1;
#10 a = 10883; b = 36285; cin = 1;
#10 a = 52325; b = 29806; cin = 1;
#10 a = 56058; b = 3454; cin = 1;
#10 a = 14236; b = 37246; cin = 0;
#10 a = 49877; b = 53281; cin = 0;
#10 a = 43754; b = 68290; cin = 0;
#10 a = 13908; b = 49088; cin = 0;
#10 a = 40389; b = 9698; cin = 1;
#10 a = 18825; b = 44842; cin = 0;
#10 a = 65015; b = 22076; cin = 0;
#10 a = 86; b = 32959; cin = 1;
#10 a = 67191; b = 61636; cin = 0;
#10 a = 28248; b = 47694; cin = 0;
#10 a = 19445; b = 61931; cin = 1;
#10 a = 55843; b = 18160; cin = 0;
#10 a = 48175; b = 38266; cin = 1;
#10 a = 19100; b = 52174; cin = 1;
#10 a = 8434; b = 22563; cin = 1;
#10 a = 51927; b = 17741; cin = 1;
#10 a = 21687; b = 12756; cin = 1;
#10 a = 60150; b = 59194; cin = 1;
#10 a = 64897; b = 56385; cin = 1;
#10 a = 5803; b = 14633; cin = 0;
#10 a = 66516; b = 10430; cin = 1;
#10 a = 827; b = 66273; cin = 1;
#10 a = 58419; b = 20801; cin = 1;
#10 a = 20654; b = 39901; cin = 1;
#10 a = 31977; b = 48335; cin = 1;
#10 a = 52998; b = 30262; cin = 0;
#10 a = 48861; b = 51949; cin = 0;
#10 a = 43153; b = 18451; cin = 0;
#10 a = 404; b = 59701; cin = 1;
#10 a = 19291; b = 41856; cin = 0;
#10 a = 15873; b = 38372; cin = 0;
#10 a = 50738; b = 15551; cin = 1;
#10 a = 57411; b = 50323; cin = 0;
#10 a = 8702; b = 47329; cin = 1;
#10 a = 12168; b = 9307; cin = 0;
#10 a = 14549; b = 38657; cin = 0;
#10 a = 34671; b = 63871; cin = 0;
#10 a = 43901; b = 37024; cin = 1;
#10 a = 42325; b = 37428; cin = 0;
#10 a = 3486; b = 56719; cin = 1;
#10 a = 49280; b = 48945; cin = 1;
#10 a = 11856; b = 29683; cin = 1;
#10 a = 40705; b = 63447; cin = 0;
#10 a = 20356; b = 48501; cin = 1;
#10 a = 39907; b = 60669; cin = 0;
#10 a = 14146; b = 51570; cin = 0;
#10 a = 64998; b = 62593; cin = 1;
#10 a = 27800; b = 12846; cin = 1;
#10 a = 55406; b = 55171; cin = 1;
#10 a = 2712; b = 58657; cin = 0;
#10 a = 61875; b = 14289; cin = 1;
#10 a = 65763; b = 26145; cin = 1;
#10 a = 15202; b = 66851; cin = 0;
#10 a = 37668; b = 63559; cin = 1;
#10 a = 61111; b = 33466; cin = 1;
#10 a = 214; b = 23964; cin = 1;
#10 a = 47974; b = 18963; cin = 1;
#10 a = 19605; b = 23115; cin = 1;
#10 a = 28260; b = 54873; cin = 1;
#10 a = 27047; b = 57586; cin = 0;
#10 a = 12553; b = 49461; cin = 0;
#10 a = 47005; b = 21576; cin = 1;
#10 a = 17492; b = 36778; cin = 0;
#10 a = 51426; b = 50798; cin = 1;
#10 a = 63861; b = 41910; cin = 0;
#10 a = 43318; b = 42124; cin = 0;
#10 a = 4346; b = 66450; cin = 1;
#10 a = 4319; b = 16055; cin = 1;
#10 a = 40786; b = 20667; cin = 0;
#10 a = 15129; b = 47714; cin = 0;
#10 a = 48130; b = 60267; cin = 0;
#10 a = 25420; b = 13624; cin = 0;
#10 a = 5207; b = 31116; cin = 1;
#10 a = 28198; b = 12542; cin = 1;
#10 a = 68395; b = 52756; cin = 1;
#10 a = 24763; b = 2426; cin = 1;
#10 a = 5096; b = 6772; cin = 1;
#10 a = 27095; b = 57443; cin = 0;
#10 a = 25858; b = 4582; cin = 1;
#10 a = 55847; b = 19711; cin = 1;
#10 a = 49773; b = 67841; cin = 1;
#10 a = 23161; b = 69613; cin = 1;
#10 a = 18126; b = 4821; cin = 0;
#10 a = 26221; b = 9371; cin = 0;
#10 a = 15114; b = 7766; cin = 0;
#10 a = 22270; b = 8882; cin = 1;
#10 a = 1549; b = 60330; cin = 1;
#10 a = 23631; b = 17425; cin = 1;
#10 a = 61767; b = 19636; cin = 1;
#10 a = 50571; b = 51835; cin = 0;
#10 a = 63440; b = 31608; cin = 0;
#10 a = 66577; b = 54770; cin = 1;
#10 a = 59691; b = 49248; cin = 0;
#10 a = 13921; b = 5469; cin = 1;
#10 a = 50693; b = 66935; cin = 0;
#10 a = 46574; b = 19205; cin = 0;
#10 a = 44881; b = 20755; cin = 0;
#10 a = 26312; b = 20738; cin = 1;
#10 a = 65187; b = 12505; cin = 1;
#10 a = 14996; b = 39428; cin = 0;
#10 a = 54517; b = 32869; cin = 1;
#10 a = 21879; b = 5798; cin = 1;
#10 a = 58854; b = 41841; cin = 1;
#10 a = 7003; b = 55762; cin = 0;
#10 a = 10874; b = 36456; cin = 1;
#10 a = 22512; b = 59382; cin = 1;
#10 a = 43032; b = 10615; cin = 0;
#10 a = 30234; b = 36927; cin = 0;
#10 a = 58510; b = 8467; cin = 1;
#10 a = 12773; b = 69815; cin = 0;
#10 a = 18872; b = 54332; cin = 1;
#10 a = 56579; b = 6211; cin = 1;
#10 a = 55408; b = 41418; cin = 1;
#10 a = 9837; b = 24773; cin = 1;
#10 a = 39735; b = 35647; cin = 1;
#10 a = 42920; b = 58160; cin = 1;
#10 a = 41663; b = 7544; cin = 0;
#10 a = 61161; b = 37779; cin = 0;
#10 a = 31397; b = 2641; cin = 1;
#10 a = 60491; b = 15414; cin = 0;
#10 a = 59013; b = 34286; cin = 1;
#10 a = 66756; b = 67217; cin = 0;
#10 a = 56649; b = 28977; cin = 0;
#10 a = 18384; b = 15166; cin = 1;
#10 a = 35882; b = 31253; cin = 1;
#10 a = 66187; b = 4174; cin = 1;
#10 a = 62227; b = 45837; cin = 1;
#10 a = 68881; b = 13351; cin = 0;
#10 a = 42463; b = 21100; cin = 1;
#10 a = 47216; b = 11591; cin = 0;
#10 a = 5433; b = 46956; cin = 0;
#10 a = 40686; b = 43712; cin = 0;
#10 a = 35798; b = 6714; cin = 1;
#10 a = 25033; b = 25098; cin = 0;
#10 a = 62688; b = 37332; cin = 1;
#10 a = 18695; b = 33520; cin = 1;
#10 a = 32862; b = 2099; cin = 1;
#10 a = 54574; b = 980; cin = 0;
#10 a = 44064; b = 19796; cin = 0;
#10 a = 36196; b = 67012; cin = 0;
#10 a = 20094; b = 48797; cin = 0;
#10 a = 14630; b = 19483; cin = 1;
#10 a = 6384; b = 31634; cin = 1;
#10 a = 3468; b = 56667; cin = 1;
#10 a = 15718; b = 25707; cin = 0;
#10 a = 59221; b = 44403; cin = 0;
#10 a = 13251; b = 7265; cin = 1;
#10 a = 59470; b = 61839; cin = 1;
#10 a = 25392; b = 12256; cin = 1;
#10 a = 36062; b = 48452; cin = 0;
#10 a = 34676; b = 44898; cin = 1;
#10 a = 56599; b = 59528; cin = 1;
#10 a = 52234; b = 42265; cin = 1;
#10 a = 54583; b = 22085; cin = 0;
#10 a = 58382; b = 14155; cin = 1;
#10 a = 29514; b = 3376; cin = 0;
#10 a = 34166; b = 62979; cin = 0;
#10 a = 17269; b = 28801; cin = 1;
#10 a = 47705; b = 54193; cin = 1;
#10 a = 27936; b = 20256; cin = 1;
#10 a = 27884; b = 31284; cin = 1;
#10 a = 6630; b = 17883; cin = 0;
#10 a = 4859; b = 46469; cin = 1;
#10 a = 57426; b = 31052; cin = 0;
#10 a = 26660; b = 65787; cin = 1;
#10 a = 67953; b = 25301; cin = 1;
#10 a = 13650; b = 35820; cin = 1;
#10 a = 59316; b = 53089; cin = 0;
#10 a = 26821; b = 7146; cin = 0;
#10 a = 52935; b = 11435; cin = 0;
#10 a = 57500; b = 39319; cin = 0;
#10 a = 59668; b = 45949; cin = 0;
#10 a = 51364; b = 27160; cin = 1;
#10 a = 15325; b = 14586; cin = 0;
#10 a = 47723; b = 41246; cin = 1;
#10 a = 628; b = 15552; cin = 0;
#10 a = 26909; b = 5554; cin = 0;
#10 a = 22522; b = 64870; cin = 0;
#10 a = 46937; b = 68043; cin = 0;
#10 a = 31897; b = 50978; cin = 1;
#10 a = 13465; b = 14831; cin = 1;
#10 a = 26317; b = 4499; cin = 0;
#10 a = 9757; b = 55863; cin = 1;
#10 a = 63315; b = 47540; cin = 1;
#10 a = 30629; b = 1615; cin = 0;
#10 a = 63730; b = 2243; cin = 0;
#10 a = 52132; b = 29152; cin = 0;
#10 a = 6355; b = 51675; cin = 0;
#10 a = 60019; b = 4964; cin = 1;
#10 a = 27181; b = 36861; cin = 0;
#10 a = 5779; b = 50326; cin = 1;
#10 a = 23696; b = 6643; cin = 0;
#10 a = 63914; b = 16401; cin = 1;
#10 a = 61293; b = 56068; cin = 1;
#10 a = 3259; b = 63049; cin = 0;
#10 a = 9175; b = 56779; cin = 1;
#10 a = 30643; b = 15263; cin = 1;
#10 a = 57665; b = 21618; cin = 0;
#10 a = 9557; b = 57989; cin = 0;
#10 a = 5844; b = 61523; cin = 1;
#10 a = 29462; b = 67302; cin = 1;
#10 a = 67911; b = 20998; cin = 1;
#10 a = 40859; b = 61264; cin = 0;
#10 a = 46022; b = 52558; cin = 0;
#10 a = 5077; b = 32169; cin = 1;
#10 a = 35747; b = 17696; cin = 0;
#10 a = 68660; b = 48339; cin = 1;
#10 a = 60726; b = 36004; cin = 0;
#10 a = 10818; b = 21913; cin = 1;
#10 a = 35875; b = 4109; cin = 0;
#10 a = 4144; b = 33572; cin = 0;
#10 a = 46388; b = 31483; cin = 0;
#10 a = 47979; b = 48695; cin = 1;
#10 a = 42323; b = 1069; cin = 1;
#10 a = 22735; b = 6147; cin = 0;
#10 a = 66196; b = 41894; cin = 0;
#10 a = 2788; b = 40555; cin = 1;
#10 a = 995; b = 7633; cin = 1;
#10 a = 44469; b = 18451; cin = 0;
#10 a = 28637; b = 30678; cin = 1;
#10 a = 4327; b = 34823; cin = 1;
#10 a = 47320; b = 57563; cin = 1;
#10 a = 17662; b = 11894; cin = 0;
#10 a = 49269; b = 54217; cin = 1;
#10 a = 39786; b = 6952; cin = 0;
#10 a = 38824; b = 49500; cin = 1;
#10 a = 55558; b = 28640; cin = 0;
#10 a = 50631; b = 29635; cin = 1;
#10 a = 34412; b = 50457; cin = 0;
#10 a = 40106; b = 55446; cin = 1;
#10 a = 49910; b = 59773; cin = 0;
#10 a = 69637; b = 37093; cin = 1;
#10 a = 27200; b = 54756; cin = 1;
#10 a = 33458; b = 10377; cin = 0;
#10 a = 17138; b = 50164; cin = 0;
#10 a = 6964; b = 65340; cin = 0;
#10 a = 38685; b = 50899; cin = 0;
#10 a = 17313; b = 7882; cin = 1;
#10 a = 3574; b = 42295; cin = 0;
#10 a = 54639; b = 58753; cin = 0;
#10 a = 66382; b = 38663; cin = 0;
#10 a = 19300; b = 14653; cin = 1;
#10 a = 6133; b = 41853; cin = 1;
#10 a = 4860; b = 51664; cin = 1;
#10 a = 57804; b = 68802; cin = 1;
#10 a = 24052; b = 5766; cin = 1;
#10 a = 39800; b = 20804; cin = 0;
#10 a = 60540; b = 38117; cin = 1;
#10 a = 17267; b = 18044; cin = 0;
#10 a = 804; b = 2683; cin = 1;
#10 a = 63434; b = 45417; cin = 1;
#10 a = 22190; b = 41069; cin = 0;
#10 a = 64392; b = 23554; cin = 1;
#10 a = 21349; b = 28414; cin = 1;
#10 a = 35036; b = 16218; cin = 1;
#10 a = 28887; b = 40270; cin = 0;
#10 a = 64431; b = 56422; cin = 0;
#10 a = 57225; b = 23314; cin = 1;
#10 a = 57902; b = 16933; cin = 1;
#10 a = 53578; b = 17737; cin = 0;
#10 a = 61656; b = 57524; cin = 1;
#10 a = 14749; b = 56066; cin = 0;
#10 a = 52495; b = 50458; cin = 0;
#10 a = 38446; b = 48160; cin = 0;
#10 a = 52414; b = 13196; cin = 0;
#10 a = 65183; b = 18436; cin = 0;
#10 a = 60071; b = 59219; cin = 0;
#10 a = 5763; b = 22796; cin = 0;
#10 a = 12277; b = 57051; cin = 0;
#10 a = 60482; b = 40629; cin = 1;
#10 a = 17723; b = 8637; cin = 1;
#10 a = 66732; b = 23386; cin = 0;
#10 a = 16811; b = 52233; cin = 0;
#10 a = 60443; b = 67032; cin = 0;
#10 a = 38842; b = 49446; cin = 1;
#10 a = 33458; b = 44629; cin = 1;
#10 a = 44697; b = 11053; cin = 0;
#10 a = 18709; b = 63168; cin = 0;
#10 a = 16036; b = 5445; cin = 1;
#10 a = 30296; b = 65928; cin = 1;
#10 a = 38645; b = 60003; cin = 0;
#10 a = 58167; b = 56735; cin = 1;
#10 a = 16459; b = 49898; cin = 0;
#10 a = 25209; b = 40342; cin = 0;
#10 a = 12120; b = 55536; cin = 0;
#10 a = 34931; b = 18994; cin = 0;
#10 a = 6178; b = 40043; cin = 1;
#10 a = 12996; b = 58753; cin = 1;
#10 a = 42610; b = 4789; cin = 1;
#10 a = 59276; b = 11437; cin = 1;
#10 a = 22923; b = 50082; cin = 0;
#10 a = 65207; b = 14601; cin = 1;
#10 a = 60878; b = 31060; cin = 0;
#10 a = 15135; b = 56270; cin = 0;
#10 a = 36423; b = 44742; cin = 0;
#10 a = 37158; b = 9673; cin = 0;
#10 a = 58874; b = 62203; cin = 0;
#10 a = 21643; b = 5199; cin = 1;
#10 a = 23932; b = 24161; cin = 0;
#10 a = 55315; b = 59789; cin = 1;
#10 a = 35330; b = 59064; cin = 1;
#10 a = 5348; b = 54272; cin = 1;
#10 a = 8454; b = 21502; cin = 1;
#10 a = 61458; b = 12989; cin = 1;
#10 a = 61156; b = 49413; cin = 1;
#10 a = 46390; b = 62923; cin = 0;
#10 a = 26970; b = 51797; cin = 1;
#10 a = 47594; b = 49792; cin = 0;
#10 a = 56971; b = 3724; cin = 0;
#10 a = 23841; b = 59040; cin = 1;
#10 a = 25796; b = 722; cin = 0;
#10 a = 54186; b = 6071; cin = 0;
#10 a = 27177; b = 14525; cin = 0;
#10 a = 7580; b = 5983; cin = 0;
#10 a = 44254; b = 43491; cin = 1;
#10 a = 32021; b = 66233; cin = 0;
#10 a = 5814; b = 69555; cin = 1;
#10 a = 41809; b = 47150; cin = 1;
#10 a = 59356; b = 10473; cin = 1;
#10 a = 7416; b = 34315; cin = 1;
#10 a = 15265; b = 36463; cin = 0;
#10 a = 58531; b = 20649; cin = 1;
#10 a = 62421; b = 24178; cin = 0;
#10 a = 17814; b = 8111; cin = 1;
#10 a = 32548; b = 28717; cin = 0;
#10 a = 3047; b = 60738; cin = 1;
#10 a = 36469; b = 42904; cin = 0;
#10 a = 51688; b = 14714; cin = 0;
#10 a = 46699; b = 50422; cin = 0;
#10 a = 45434; b = 57838; cin = 1;
#10 a = 9562; b = 49455; cin = 0;
#10 a = 44412; b = 14339; cin = 0;
#10 a = 61685; b = 6760; cin = 0;
#10 a = 47131; b = 926; cin = 1;
#10 a = 61264; b = 9826; cin = 0;
#10 a = 2536; b = 12873; cin = 1;
#10 a = 56393; b = 49342; cin = 1;
#10 a = 39805; b = 31030; cin = 1;
#10 a = 46720; b = 54081; cin = 1;
#10 a = 64108; b = 29516; cin = 1;
#10 a = 22163; b = 15430; cin = 1;
#10 a = 63033; b = 36194; cin = 0;
#10 a = 54553; b = 27879; cin = 0;
#10 a = 46604; b = 51362; cin = 1;
#10 a = 46765; b = 42626; cin = 1;
#10 a = 5644; b = 21514; cin = 1;
#10 a = 25261; b = 7907; cin = 1;
#10 a = 64134; b = 24064; cin = 0;
#10 a = 24074; b = 784; cin = 1;
#10 a = 58083; b = 41244; cin = 1;
#10 a = 32635; b = 39759; cin = 1;
#10 a = 32994; b = 32793; cin = 1;
#10 a = 1340; b = 17346; cin = 0;
#10 a = 69150; b = 63950; cin = 0;
#10 a = 67887; b = 40716; cin = 0;
#10 a = 6451; b = 46360; cin = 0;
#10 a = 4240; b = 47973; cin = 1;
#10 a = 51371; b = 18459; cin = 0;
#10 a = 35885; b = 42533; cin = 0;
#10 a = 50833; b = 6969; cin = 1;
#10 a = 1648; b = 15956; cin = 0;
#10 a = 37894; b = 48950; cin = 1;
#10 a = 16685; b = 26642; cin = 0;
#10 a = 23356; b = 25792; cin = 0;
#10 a = 11388; b = 23680; cin = 0;
#10 a = 18399; b = 6483; cin = 0;
#10 a = 46923; b = 10723; cin = 1;
#10 a = 59707; b = 62094; cin = 1;
#10 a = 2907; b = 4332; cin = 0;
#10 a = 16891; b = 31517; cin = 1;
#10 a = 48472; b = 33165; cin = 1;
#10 a = 26165; b = 1059; cin = 1;
#10 a = 36650; b = 17745; cin = 1;
#10 a = 64482; b = 17453; cin = 0;
#10 a = 62617; b = 28841; cin = 0;
#10 a = 7819; b = 23592; cin = 1;
#10 a = 45734; b = 46868; cin = 0;
#10 a = 37973; b = 12927; cin = 0;
#10 a = 48672; b = 15834; cin = 0;
#10 a = 31905; b = 9077; cin = 1;
#10 a = 68458; b = 33902; cin = 1;
#10 a = 50968; b = 60067; cin = 0;
#10 a = 12427; b = 26717; cin = 1;
#10 a = 529; b = 21200; cin = 0;
#10 a = 14423; b = 60169; cin = 0;
#10 a = 28349; b = 44340; cin = 0;
#10 a = 25110; b = 66426; cin = 0;
#10 a = 56242; b = 10752; cin = 1;
#10 a = 32172; b = 59424; cin = 1;
#10 a = 12435; b = 67681; cin = 1;
#10 a = 566; b = 42492; cin = 1;
#10 a = 21863; b = 23460; cin = 0;
#10 a = 44220; b = 35887; cin = 1;
#10 a = 37025; b = 36416; cin = 1;
#10 a = 932; b = 27191; cin = 0;
#10 a = 40032; b = 31892; cin = 1;
#10 a = 9076; b = 57002; cin = 1;
#10 a = 1341; b = 19596; cin = 1;
#10 a = 6532; b = 51769; cin = 0;
#10 a = 3910; b = 64204; cin = 1;
#10 a = 10365; b = 64770; cin = 1;
#10 a = 50722; b = 62986; cin = 1;
#10 a = 57498; b = 13558; cin = 1;
#10 a = 44639; b = 50583; cin = 1;
#10 a = 5685; b = 27867; cin = 1;
#10 a = 50547; b = 67899; cin = 1;
#10 a = 22454; b = 53328; cin = 0;
#10 a = 14436; b = 31021; cin = 0;
#10 a = 63521; b = 37553; cin = 1;
#10 a = 32031; b = 17815; cin = 1;
#10 a = 44575; b = 4532; cin = 0;
#10 a = 29610; b = 31606; cin = 0;
#10 a = 14458; b = 19104; cin = 0;
#10 a = 35193; b = 40096; cin = 1;
#10 a = 68696; b = 45781; cin = 1;
#10 a = 35743; b = 2680; cin = 0;
#10 a = 34683; b = 25135; cin = 0;
#10 a = 66977; b = 15923; cin = 1;
#10 a = 48867; b = 9444; cin = 1;
#10 a = 36175; b = 17828; cin = 0;
#10 a = 40390; b = 38755; cin = 1;
#10 a = 39376; b = 68365; cin = 1;
#10 a = 7700; b = 59175; cin = 0;
#10 a = 59582; b = 24368; cin = 0;
#10 a = 22048; b = 69417; cin = 1;
#10 a = 58733; b = 11512; cin = 1;
#10 a = 23317; b = 22547; cin = 0;
#10 a = 17582; b = 19524; cin = 1;
#10 a = 42867; b = 68392; cin = 0;
#10 a = 12058; b = 10919; cin = 0;
#10 a = 45417; b = 27661; cin = 1;
#10 a = 13308; b = 43390; cin = 0;
#10 a = 12805; b = 51090; cin = 0;
#10 a = 31407; b = 17025; cin = 0;
#10 a = 66457; b = 39073; cin = 1;
#10 a = 30936; b = 4158; cin = 0;
#10 a = 44448; b = 27475; cin = 1;
#10 a = 13094; b = 45057; cin = 0;
#10 a = 44016; b = 64277; cin = 0;
#10 a = 38030; b = 6335; cin = 1;
#10 a = 2576; b = 51752; cin = 0;
#10 a = 29525; b = 41412; cin = 0;
#10 a = 31191; b = 54218; cin = 1;
#10 a = 68385; b = 61977; cin = 0;
#10 a = 59948; b = 58435; cin = 1;
#10 a = 3631; b = 65723; cin = 1;
#10 a = 28827; b = 40171; cin = 0;
#10 a = 6571; b = 29618; cin = 0;
#10 a = 50191; b = 3634; cin = 1;
#10 a = 22203; b = 18016; cin = 0;
#10 a = 27838; b = 20592; cin = 1;
#10 a = 61134; b = 26469; cin = 1;
#10 a = 21469; b = 34012; cin = 1;
#10 a = 55598; b = 32398; cin = 1;
#10 a = 60400; b = 68698; cin = 0;
#10 a = 56979; b = 2329; cin = 1;
#10 a = 11364; b = 31157; cin = 1;
#10 a = 39576; b = 37728; cin = 1;
#10 a = 19198; b = 17919; cin = 1;
#10 a = 63097; b = 16474; cin = 1;
#10 a = 43332; b = 20664; cin = 1;
#10 a = 51671; b = 11798; cin = 0;
#10 a = 31422; b = 9619; cin = 0;
#10 a = 41744; b = 65217; cin = 0;
#10 a = 44043; b = 31969; cin = 0;
#10 a = 34777; b = 18948; cin = 0;
#10 a = 21234; b = 6664; cin = 1;
#10 a = 567; b = 22593; cin = 1;
#10 a = 9518; b = 41791; cin = 0;
#10 a = 68455; b = 34889; cin = 0;
#10 a = 5408; b = 54573; cin = 0;
#10 a = 55657; b = 36244; cin = 0;
#10 a = 62375; b = 44018; cin = 0;
#10 a = 56754; b = 62114; cin = 1;
#10 a = 36234; b = 12509; cin = 1;
#10 a = 38061; b = 47286; cin = 1;
#10 a = 18569; b = 44873; cin = 0;
#10 a = 6586; b = 45440; cin = 1;
#10 a = 8683; b = 31311; cin = 0;
#10 a = 28699; b = 29766; cin = 1;
#10 a = 17893; b = 35175; cin = 0;
#10 a = 27751; b = 67184; cin = 0;
#10 a = 49407; b = 59560; cin = 1;
#10 a = 10683; b = 22666; cin = 1;
#10 a = 37177; b = 58900; cin = 1;
#10 a = 1992; b = 3313; cin = 1;
#10 a = 9403; b = 68234; cin = 0;
#10 a = 69831; b = 4820; cin = 1;
#10 a = 59204; b = 59855; cin = 0;
#10 a = 44017; b = 64906; cin = 0;
#10 a = 16422; b = 12799; cin = 1;
#10 a = 43401; b = 40550; cin = 0;
#10 a = 12975; b = 19958; cin = 0;
#10 a = 2920; b = 30641; cin = 0;
#10 a = 31332; b = 44170; cin = 0;
#10 a = 25901; b = 46162; cin = 0;
#10 a = 20460; b = 31918; cin = 0;
#10 a = 59893; b = 8101; cin = 1;
#10 a = 27470; b = 67306; cin = 0;
#10 a = 50006; b = 17675; cin = 1;
#10 a = 8660; b = 34097; cin = 0;
#10 a = 2490; b = 53850; cin = 1;
#10 a = 39856; b = 43178; cin = 1;
#10 a = 66782; b = 46098; cin = 0;
#10 a = 22726; b = 7430; cin = 1;
#10 a = 37570; b = 9683; cin = 1;
#10 a = 55728; b = 6496; cin = 1;
#10 a = 48473; b = 42741; cin = 1;
#10 a = 22390; b = 211; cin = 1;
#10 a = 9810; b = 50217; cin = 0;
#10 a = 38489; b = 58877; cin = 1;
#10 a = 9968; b = 37719; cin = 0;
#10 a = 68349; b = 7575; cin = 0;
#10 a = 6688; b = 50709; cin = 0;
#10 a = 22020; b = 3435; cin = 1;
#10 a = 11523; b = 41006; cin = 0;
#10 a = 47189; b = 3086; cin = 0;
#10 a = 21124; b = 27911; cin = 1;
#10 a = 49513; b = 50301; cin = 0;
#10 a = 5208; b = 36464; cin = 1;
#10 a = 48578; b = 4953; cin = 1;
#10 a = 32398; b = 61273; cin = 0;
#10 a = 68; b = 59622; cin = 0;
#10 a = 57268; b = 66310; cin = 1;
#10 a = 20566; b = 18331; cin = 1;
#10 a = 37647; b = 29854; cin = 1;
#10 a = 17116; b = 53395; cin = 1;
#10 a = 26728; b = 50872; cin = 1;
#10 a = 55434; b = 30385; cin = 0;
#10 a = 37998; b = 11946; cin = 0;
#10 a = 23484; b = 60524; cin = 0;
#10 a = 67847; b = 22922; cin = 1;
#10 a = 56281; b = 69342; cin = 0;
#10 a = 28643; b = 56610; cin = 0;
#10 a = 51715; b = 53529; cin = 1;
#10 a = 54574; b = 67528; cin = 0;
#10 a = 28439; b = 14644; cin = 1;
#10 a = 51742; b = 41373; cin = 1;
#10 a = 9309; b = 26807; cin = 1;
#10 a = 63530; b = 41157; cin = 1;
#10 a = 37862; b = 40993; cin = 1;
#10 a = 63500; b = 15192; cin = 0;
#10 a = 56764; b = 47826; cin = 0;
#10 a = 63298; b = 6469; cin = 1;
#10 a = 18846; b = 34536; cin = 0;
#10 a = 62726; b = 19110; cin = 0;
#10 a = 42812; b = 47549; cin = 1;
#10 a = 52645; b = 5644; cin = 0;
#10 a = 43351; b = 61305; cin = 1;
#10 a = 40794; b = 54835; cin = 0;
#10 a = 26535; b = 69050; cin = 0;
#10 a = 26448; b = 62550; cin = 0;
#10 a = 25636; b = 25666; cin = 0;
#10 a = 519; b = 65316; cin = 0;
#10 a = 32012; b = 14163; cin = 0;
#10 a = 47034; b = 53241; cin = 1;
#10 a = 35936; b = 26053; cin = 0;
#10 a = 63131; b = 55050; cin = 0;
#10 a = 14403; b = 28401; cin = 0;
#10 a = 38834; b = 45547; cin = 1;
#10 a = 34423; b = 48434; cin = 1;
#10 a = 47357; b = 4883; cin = 0;
#10 a = 51835; b = 6871; cin = 0;
#10 a = 34140; b = 7390; cin = 1;
#10 a = 22914; b = 15754; cin = 0;
#10 a = 22576; b = 39140; cin = 1;
#10 a = 41349; b = 5077; cin = 0;
#10 a = 14024; b = 44560; cin = 0;
#10 a = 38694; b = 58964; cin = 0;
#10 a = 31022; b = 27798; cin = 1;
#10 a = 8186; b = 38573; cin = 0;
#10 a = 54399; b = 15930; cin = 1;
#10 a = 45867; b = 44118; cin = 0;
#10 a = 16650; b = 8258; cin = 1;
#10 a = 29101; b = 31172; cin = 1;
#10 a = 55715; b = 30100; cin = 0;
#10 a = 65570; b = 47802; cin = 1;
#10 a = 7830; b = 61826; cin = 1;
#10 a = 5140; b = 6872; cin = 1;
#10 a = 7204; b = 37895; cin = 0;
#10 a = 31168; b = 46081; cin = 1;
#10 a = 33566; b = 6832; cin = 0;
#10 a = 40847; b = 29052; cin = 0;
#10 a = 7703; b = 45702; cin = 0;
#10 a = 51950; b = 51155; cin = 0;
#10 a = 18304; b = 36870; cin = 0;
#10 a = 23798; b = 8792; cin = 0;
#10 a = 34369; b = 16622; cin = 0;
#10 a = 19500; b = 68114; cin = 1;
#10 a = 39948; b = 5319; cin = 0;
#10 a = 18194; b = 36487; cin = 1;
#10 a = 35013; b = 53; cin = 1;
#10 a = 44115; b = 17252; cin = 1;
#10 a = 3687; b = 24955; cin = 1;
#10 a = 65165; b = 53258; cin = 0;
#10 a = 40519; b = 47914; cin = 0;
#10 a = 45974; b = 1712; cin = 0;
#10 a = 29230; b = 36081; cin = 0;
#10 a = 50665; b = 31933; cin = 1;
#10 a = 55324; b = 1881; cin = 0;
#10 a = 27878; b = 20075; cin = 1;
#10 a = 22865; b = 31441; cin = 0;
#10 a = 1036; b = 5556; cin = 0;
#10 a = 8260; b = 55596; cin = 1;
#10 a = 61185; b = 27113; cin = 1;
#10 a = 1618; b = 67633; cin = 1;
#10 a = 25272; b = 19959; cin = 1;
#10 a = 57719; b = 25541; cin = 0;
#10 a = 13139; b = 6206; cin = 0;
#10 a = 13026; b = 37882; cin = 1;
#10 a = 18232; b = 65760; cin = 1;
#10 a = 36277; b = 64977; cin = 0;
#10 a = 54375; b = 66014; cin = 0;
#10 a = 42429; b = 4274; cin = 0;
#10 a = 55439; b = 41811; cin = 0;
#10 a = 28058; b = 19781; cin = 1;
#10 a = 48592; b = 45054; cin = 0;
#10 a = 47189; b = 9125; cin = 1;
#10 a = 11868; b = 68616; cin = 0;
#10 a = 8480; b = 11643; cin = 0;
#10 a = 53325; b = 6227; cin = 1;
#10 a = 48246; b = 42505; cin = 0;
#10 a = 50960; b = 3232; cin = 0;
#10 a = 59231; b = 45662; cin = 0;
#10 a = 53097; b = 31101; cin = 0;
#10 a = 50429; b = 35511; cin = 1;
#10 a = 21746; b = 14103; cin = 1;
#10 a = 13022; b = 61293; cin = 0;
#10 a = 29840; b = 49513; cin = 1;
#10 a = 52864; b = 34345; cin = 0;
#10 a = 20122; b = 17670; cin = 1;
#10 a = 29493; b = 42269; cin = 0;
#10 a = 33842; b = 23229; cin = 1;
#10 a = 34204; b = 12460; cin = 1;
#10 a = 15193; b = 41910; cin = 0;
#10 a = 37993; b = 68691; cin = 1;
#10 a = 56926; b = 20438; cin = 1;
#10 a = 50914; b = 33460; cin = 0;
#10 a = 30378; b = 63300; cin = 1;
#10 a = 54811; b = 22516; cin = 0;
#10 a = 67239; b = 18991; cin = 0;
#10 a = 39543; b = 48484; cin = 1;
#10 a = 30703; b = 58678; cin = 1;
#10 a = 1448; b = 22883; cin = 1;
#10 a = 41503; b = 38076; cin = 1;
#10 a = 19011; b = 52421; cin = 1;
#10 a = 32031; b = 39347; cin = 1;
#10 a = 35506; b = 66613; cin = 1;
#10 a = 30274; b = 3344; cin = 0;
#10 a = 50907; b = 58155; cin = 0;
#10 a = 35885; b = 55395; cin = 1;
#10 a = 38533; b = 1290; cin = 0;
#10 a = 59803; b = 8345; cin = 0;
#10 a = 10654; b = 9794; cin = 1;
#10 a = 20317; b = 27649; cin = 1;
#10 a = 1891; b = 46661; cin = 0;
#10 a = 28508; b = 55044; cin = 0;
#10 a = 29211; b = 20550; cin = 1;
#10 a = 16078; b = 27176; cin = 1;
#10 a = 19894; b = 54435; cin = 1;
#10 a = 22579; b = 20320; cin = 0;
#10 a = 44254; b = 58853; cin = 0;
#10 a = 20766; b = 25008; cin = 1;
#10 a = 55957; b = 12014; cin = 1;
#10 a = 20382; b = 32332; cin = 1;
#10 a = 22884; b = 10575; cin = 0;
#10 a = 30510; b = 39083; cin = 0;
#10 a = 7484; b = 44646; cin = 0;
#10 a = 51072; b = 60724; cin = 0;
#10 a = 4355; b = 10619; cin = 1;
#10 a = 15794; b = 33198; cin = 1;
#10 a = 58980; b = 53804; cin = 0;
#10 a = 56160; b = 4571; cin = 1;
#10 a = 61686; b = 60528; cin = 1;
#10 a = 53357; b = 10910; cin = 1;
#10 a = 2678; b = 10146; cin = 0;
#10 a = 45012; b = 17009; cin = 1;
#10 a = 48742; b = 24493; cin = 1;
#10 a = 3022; b = 5565; cin = 0;
#10 a = 30830; b = 9921; cin = 1;
#10 a = 43073; b = 2067; cin = 1;
#10 a = 51988; b = 37400; cin = 1;
#10 a = 49757; b = 23560; cin = 0;
#10 a = 48886; b = 15246; cin = 0;
#10 a = 13677; b = 68604; cin = 1;
#10 a = 57153; b = 1282; cin = 1;
#10 a = 41203; b = 22647; cin = 0;
#10 a = 40689; b = 1389; cin = 0;
#10 a = 38468; b = 4412; cin = 1;
#10 a = 3324; b = 11594; cin = 0;
#10 a = 25151; b = 31020; cin = 0;
#10 a = 10176; b = 13008; cin = 0;
#10 a = 25358; b = 62765; cin = 0;
#10 a = 68758; b = 41651; cin = 1;
#10 a = 55391; b = 31681; cin = 1;
#10 a = 52934; b = 65186; cin = 1;
#10 a = 36975; b = 12741; cin = 0;
#10 a = 38026; b = 53430; cin = 0;
#10 a = 39922; b = 68251; cin = 0;
#10 a = 47383; b = 47927; cin = 0;
#10 a = 64766; b = 3079; cin = 0;
#10 a = 36920; b = 59607; cin = 1;
#10 a = 122; b = 14965; cin = 0;
#10 a = 56884; b = 60076; cin = 0;
#10 a = 35245; b = 45467; cin = 1;
#10 a = 12210; b = 4753; cin = 1;
#10 a = 36810; b = 18080; cin = 0;
#10 a = 60408; b = 56106; cin = 1;
#10 a = 15396; b = 2380; cin = 0;
#10 a = 44796; b = 49764; cin = 1;
#10 a = 62143; b = 20882; cin = 0;
#10 a = 40509; b = 57802; cin = 0;
#10 a = 8236; b = 57924; cin = 1;
#10 a = 38729; b = 21160; cin = 1;
#10 a = 17225; b = 32758; cin = 0;
#10 a = 27402; b = 21320; cin = 1;
#10 a = 55469; b = 34482; cin = 0;
#10 a = 26277; b = 24891; cin = 0;
#10 a = 50516; b = 40287; cin = 1;
#10 a = 25710; b = 61436; cin = 1;
#10 a = 2480; b = 29931; cin = 1;
#10 a = 5032; b = 440; cin = 1;
#10 a = 67192; b = 55029; cin = 1;
#10 a = 4318; b = 23758; cin = 1;
#10 a = 1519; b = 40983; cin = 1;
#10 a = 66892; b = 44737; cin = 0;
#10 a = 67017; b = 30206; cin = 0;
#10 a = 15223; b = 32835; cin = 1;
#10 a = 65888; b = 13352; cin = 1;
#10 a = 48933; b = 39062; cin = 1;
#10 a = 11742; b = 17894; cin = 0;
#10 a = 65433; b = 22927; cin = 0;
#10 a = 13278; b = 20119; cin = 1;
#10 a = 65399; b = 789; cin = 1;
#10 a = 68680; b = 48661; cin = 0;
#10 a = 34720; b = 45553; cin = 1;
#10 a = 68432; b = 42570; cin = 1;
#10 a = 66626; b = 57794; cin = 1;
#10 a = 43360; b = 53682; cin = 1;
#10 a = 13085; b = 32615; cin = 1;
#10 a = 44246; b = 20709; cin = 0;
#10 a = 35338; b = 62494; cin = 1;
#10 a = 26870; b = 5772; cin = 0;
#10 a = 49784; b = 47523; cin = 0;
#10 a = 2807; b = 46203; cin = 1;
#10 a = 66814; b = 57275; cin = 0;
#10 a = 11909; b = 32059; cin = 0;
#10 a = 33563; b = 28686; cin = 0;
#10 a = 18052; b = 48398; cin = 0;
#10 a = 15893; b = 61483; cin = 1;
#10 a = 5500; b = 35729; cin = 0;
#10 a = 13002; b = 1067; cin = 0;
#10 a = 19783; b = 4289; cin = 0;
#10 a = 23036; b = 30425; cin = 1;
#10 a = 27078; b = 9585; cin = 1;
#10 a = 9781; b = 6399; cin = 0;
#10 a = 38037; b = 64660; cin = 0;
#10 a = 15215; b = 28223; cin = 0;
#10 a = 50188; b = 46275; cin = 0;
#10 a = 45194; b = 38520; cin = 1;
#10 a = 49168; b = 44021; cin = 0;
#10 a = 50202; b = 33375; cin = 1;
#10 a = 67379; b = 29511; cin = 0;
#10 a = 43031; b = 52547; cin = 0;
#10 a = 19855; b = 9625; cin = 1;
#10 a = 65586; b = 65758; cin = 0;
#10 a = 28592; b = 33795; cin = 0;
#10 a = 23658; b = 49010; cin = 0;
#10 a = 23762; b = 5550; cin = 1;
#10 a = 25912; b = 50745; cin = 0;
#10 a = 65897; b = 6265; cin = 1;
#10 a = 47963; b = 56467; cin = 0;
#10 a = 7448; b = 30198; cin = 1;
#10 a = 17575; b = 3230; cin = 0;
#10 a = 58127; b = 69437; cin = 1;
#10 a = 38264; b = 65023; cin = 1;
#10 a = 1152; b = 69967; cin = 0;
#10 a = 28700; b = 69978; cin = 1;
#10 a = 60824; b = 23740; cin = 1;
#10 a = 22872; b = 26005; cin = 0;
#10 a = 46144; b = 68254; cin = 1;
#10 a = 43437; b = 22570; cin = 1;
#10 a = 50457; b = 30018; cin = 1;
#10 a = 16989; b = 47593; cin = 1;
#10 a = 36067; b = 12072; cin = 0;
#10 a = 17475; b = 26688; cin = 1;
#10 a = 64640; b = 4192; cin = 1;
#10 a = 5601; b = 32893; cin = 1;
#10 a = 41924; b = 69; cin = 1;
#10 a = 60149; b = 22941; cin = 0;
#10 a = 59120; b = 45437; cin = 1;
#10 a = 64355; b = 18874; cin = 1;
#10 a = 8762; b = 69332; cin = 1;
#10 a = 7016; b = 16321; cin = 1;
#10 a = 31203; b = 28740; cin = 1;
#10 a = 54828; b = 22567; cin = 0;
#10 a = 3475; b = 63560; cin = 0;
#10 a = 44794; b = 45513; cin = 1;
#10 a = 39739; b = 63789; cin = 1;
#10 a = 34777; b = 53938; cin = 0;
#10 a = 32171; b = 43058; cin = 0;
#10 a = 4172; b = 37414; cin = 0;
#10 a = 22391; b = 46176; cin = 0;
#10 a = 23333; b = 29544; cin = 1;
#10 a = 48220; b = 37100; cin = 0;
#10 a = 15179; b = 21928; cin = 1;
#10 a = 8827; b = 1755; cin = 1;
#10 a = 6668; b = 46550; cin = 0;
#10 a = 13753; b = 62641; cin = 1;
#10 a = 20908; b = 3770; cin = 0;
#10 a = 27357; b = 35942; cin = 0;
#10 a = 55595; b = 40114; cin = 0;
#10 a = 56355; b = 38858; cin = 1;
#10 a = 9152; b = 38543; cin = 1;
#10 a = 48269; b = 16763; cin = 1;
#10 a = 46127; b = 31942; cin = 1;
#10 a = 19257; b = 40770; cin = 1;
#10 a = 9594; b = 47438; cin = 1;
#10 a = 21797; b = 37543; cin = 0;
#10 a = 27788; b = 34804; cin = 1;
#10 a = 17718; b = 38513; cin = 1;
#10 a = 50707; b = 24108; cin = 1;
#10 a = 51109; b = 10463; cin = 1;
#10 a = 50392; b = 19615; cin = 0;
#10 a = 9220; b = 44237; cin = 1;
#10 a = 51499; b = 66716; cin = 0;
#10 a = 45707; b = 15973; cin = 0;
#10 a = 18022; b = 1920; cin = 0;
#10 a = 36887; b = 23717; cin = 1;
#10 a = 48393; b = 27857; cin = 1;
#10 a = 63670; b = 45576; cin = 0;
#10 a = 21241; b = 26283; cin = 0;
#10 a = 65279; b = 53744; cin = 0;
#10 a = 54526; b = 34137; cin = 1;
#10 a = 12317; b = 19709; cin = 0;
#10 a = 56870; b = 1208; cin = 1;
#10 a = 63366; b = 23267; cin = 0;
#10 a = 16984; b = 41289; cin = 0;
#10 a = 64392; b = 54528; cin = 1;
#10 a = 9344; b = 32922; cin = 1;
#10 a = 35451; b = 2944; cin = 1;
#10 a = 53720; b = 24186; cin = 0;
#10 a = 2448; b = 65817; cin = 0;
#10 a = 7992; b = 50343; cin = 1;
#10 a = 9504; b = 39012; cin = 0;
#10 a = 8900; b = 25883; cin = 1;
#10 a = 51365; b = 65601; cin = 0;
#10 a = 39804; b = 12586; cin = 0;
#10 a = 6514; b = 53330; cin = 0;
#10 a = 66942; b = 62674; cin = 0;
#10 a = 15227; b = 4478; cin = 1;
#10 a = 9088; b = 34550; cin = 1;
#10 a = 29232; b = 36998; cin = 0;
#10 a = 9472; b = 44991; cin = 1;
#10 a = 23850; b = 54495; cin = 0;
#10 a = 34288; b = 39747; cin = 1;
#10 a = 45935; b = 67465; cin = 0;
#10 a = 57202; b = 13621; cin = 0;
#10 a = 16110; b = 20135; cin = 1;
#10 a = 29546; b = 17077; cin = 1;
#10 a = 52257; b = 32304; cin = 1;
#10 a = 7912; b = 41392; cin = 1;
#10 a = 34105; b = 46976; cin = 0;
#10 a = 56115; b = 56449; cin = 1;
#10 a = 34820; b = 56651; cin = 0;
#10 a = 52538; b = 20939; cin = 1;
#10 a = 2491; b = 43227; cin = 0;
#10 a = 18046; b = 30429; cin = 1;
#10 a = 22538; b = 22891; cin = 1;
#10 a = 10361; b = 28789; cin = 0;
#10 a = 13563; b = 57398; cin = 1;
#10 a = 44890; b = 65310; cin = 1;
#10 a = 40768; b = 29415; cin = 0;
#10 a = 49996; b = 61882; cin = 1;
#10 a = 10567; b = 3055; cin = 0;
#10 a = 1985; b = 55593; cin = 1;
#10 a = 9502; b = 34437; cin = 0;
#10 a = 14485; b = 28835; cin = 1;
#10 a = 9440; b = 27725; cin = 0;
#10 a = 48179; b = 14439; cin = 0;
#10 a = 10348; b = 28002; cin = 0;
#10 a = 4821; b = 2892; cin = 1;
#10 a = 40686; b = 20012; cin = 0;
#10 a = 29880; b = 46360; cin = 1;
#10 a = 5523; b = 33279; cin = 0;
#10 a = 14169; b = 11616; cin = 1;
#10 a = 67403; b = 21119; cin = 0;
#10 a = 215; b = 11956; cin = 1;
#10 a = 9809; b = 21396; cin = 1;
#10 a = 42293; b = 45928; cin = 0;
#10 a = 9919; b = 56276; cin = 0;
#10 a = 34944; b = 61097; cin = 0;
#10 a = 31631; b = 8135; cin = 1;
#10 a = 34085; b = 38016; cin = 1;
#10 a = 28422; b = 19891; cin = 1;
#10 a = 25814; b = 34061; cin = 1;
#10 a = 55152; b = 7816; cin = 0;
#10 a = 48926; b = 8031; cin = 0;
#10 a = 47888; b = 64192; cin = 1;
#10 a = 50927; b = 12838; cin = 1;
#10 a = 22053; b = 69109; cin = 1;
#10 a = 67533; b = 10405; cin = 0;
#10 a = 22257; b = 42036; cin = 1;
#10 a = 66994; b = 52474; cin = 1;
#10 a = 64444; b = 10896; cin = 1;
#10 a = 25173; b = 36711; cin = 0;
#10 a = 67518; b = 21863; cin = 0;
#10 a = 37335; b = 47141; cin = 1;
#10 a = 65459; b = 1381; cin = 0;
#10 a = 44980; b = 52308; cin = 0;
#10 a = 46781; b = 50713; cin = 1;
#10 a = 11210; b = 48246; cin = 1;
#10 a = 36736; b = 46856; cin = 1;
#10 a = 398; b = 43850; cin = 1;
#10 a = 48427; b = 38294; cin = 0;
#10 a = 22700; b = 39819; cin = 1;
#10 a = 54682; b = 37338; cin = 0;
#10 a = 832; b = 51025; cin = 1;
#10 a = 1366; b = 22836; cin = 1;
#10 a = 66092; b = 44169; cin = 1;
#10 a = 50008; b = 20950; cin = 1;
#10 a = 33033; b = 32161; cin = 1;
#10 a = 2816; b = 68897; cin = 1;
#10 a = 60988; b = 45647; cin = 0;
#10 a = 55281; b = 427; cin = 0;
#10 a = 13175; b = 69479; cin = 0;
#10 a = 31428; b = 54162; cin = 0;
#10 a = 24248; b = 31346; cin = 1;
#10 a = 64210; b = 32712; cin = 1;
#10 a = 35553; b = 5156; cin = 0;
#10 a = 11908; b = 55164; cin = 1;
#10 a = 62625; b = 64550; cin = 0;
#10 a = 44293; b = 67366; cin = 1;
#10 a = 26464; b = 58354; cin = 1;
#10 a = 28838; b = 19988; cin = 0;
#10 a = 45859; b = 9515; cin = 1;
#10 a = 32699; b = 40944; cin = 1;
#10 a = 56877; b = 41544; cin = 0;
#10 a = 38432; b = 35754; cin = 0;
#10 a = 19175; b = 47659; cin = 1;
#10 a = 67736; b = 59568; cin = 1;
#10 a = 19951; b = 28545; cin = 1;
#10 a = 4327; b = 2838; cin = 0;
#10 a = 33952; b = 5655; cin = 0;
#10 a = 15577; b = 10845; cin = 0;
#10 a = 43981; b = 56704; cin = 0;
#10 a = 25513; b = 65755; cin = 0;
#10 a = 13910; b = 52632; cin = 0;
#10 a = 33654; b = 67416; cin = 1;
#10 a = 62463; b = 62944; cin = 0;
#10 a = 2780; b = 37032; cin = 0;
#10 a = 68261; b = 56983; cin = 0;
#10 a = 58293; b = 61310; cin = 0;
#10 a = 68395; b = 1614; cin = 1;
#10 a = 66851; b = 17192; cin = 1;
#10 a = 38000; b = 61173; cin = 1;
#10 a = 42312; b = 63038; cin = 1;
#10 a = 63920; b = 53301; cin = 1;
#10 a = 33424; b = 16955; cin = 0;
#10 a = 38683; b = 55770; cin = 0;
#10 a = 21602; b = 58550; cin = 0;
#10 a = 16792; b = 33164; cin = 1;
#10 a = 40528; b = 21457; cin = 1;
#10 a = 43455; b = 66204; cin = 1;
#10 a = 28388; b = 63055; cin = 1;
#10 a = 24167; b = 7407; cin = 1;
#10 a = 29355; b = 49719; cin = 1;
#10 a = 53946; b = 19991; cin = 0;
#10 a = 13873; b = 53416; cin = 0;
#10 a = 41217; b = 22099; cin = 0;
#10 a = 37857; b = 20053; cin = 1;
#10 a = 25177; b = 36846; cin = 1;
#10 a = 45832; b = 7374; cin = 0;
#10 a = 34149; b = 50829; cin = 0;
#10 a = 24081; b = 55570; cin = 1;
#10 a = 31204; b = 9737; cin = 1;
#10 a = 52205; b = 39092; cin = 0;
#10 a = 66245; b = 69390; cin = 0;
#10 a = 63585; b = 13264; cin = 0;
#10 a = 7881; b = 30833; cin = 1;
#10 a = 30652; b = 68691; cin = 1;
#10 a = 41973; b = 220; cin = 1;
#10 a = 16458; b = 46053; cin = 1;
#10 a = 35104; b = 56554; cin = 1;
#10 a = 3602; b = 10635; cin = 1;
#10 a = 57859; b = 18192; cin = 0;
#10 a = 3172; b = 397; cin = 1;
#10 a = 44557; b = 66642; cin = 1;
#10 a = 12285; b = 60228; cin = 1;
#10 a = 33429; b = 44461; cin = 1;
#10 a = 6672; b = 5113; cin = 0;
#10 a = 46321; b = 23438; cin = 0;
#10 a = 29168; b = 39896; cin = 1;
#10 a = 43038; b = 51352; cin = 0;
#10 a = 60441; b = 54954; cin = 1;
#10 a = 63414; b = 42814; cin = 1;
#10 a = 52476; b = 22338; cin = 1;
#10 a = 56983; b = 43247; cin = 1;
#10 a = 60881; b = 55532; cin = 1;
#10 a = 8042; b = 65313; cin = 1;
#10 a = 32389; b = 48338; cin = 0;
#10 a = 55427; b = 24659; cin = 1;
#10 a = 8686; b = 30180; cin = 1;
#10 a = 54349; b = 3218; cin = 0;
#10 a = 62919; b = 40011; cin = 0;
#10 a = 35773; b = 9777; cin = 0;
#10 a = 3170; b = 38605; cin = 1;
#10 a = 64613; b = 25589; cin = 0;
#10 a = 29051; b = 62822; cin = 1;
#10 a = 53716; b = 47216; cin = 0;
#10 a = 52843; b = 55958; cin = 0;
#10 a = 57084; b = 41385; cin = 0;
#10 a = 14763; b = 26423; cin = 0;
#10 a = 58690; b = 57125; cin = 0;
#10 a = 60322; b = 50044; cin = 1;
#10 a = 46909; b = 15817; cin = 0;
#10 a = 52661; b = 65340; cin = 1;
#10 a = 10752; b = 36305; cin = 0;
#10 a = 58443; b = 65356; cin = 0;
#10 a = 68018; b = 49073; cin = 1;
#10 a = 2906; b = 31916; cin = 1;
#10 a = 32485; b = 65352; cin = 0;
#10 a = 16723; b = 10115; cin = 0;
#10 a = 31141; b = 45158; cin = 1;
#10 a = 1481; b = 35480; cin = 1;
#10 a = 11832; b = 12389; cin = 1;
#10 a = 8312; b = 65051; cin = 1;
#10 a = 43397; b = 5803; cin = 0;
#10 a = 56776; b = 40598; cin = 1;
#10 a = 62976; b = 38616; cin = 0;
#10 a = 46393; b = 17875; cin = 0;
#10 a = 62120; b = 50360; cin = 1;
#10 a = 49233; b = 67083; cin = 0;
#10 a = 62769; b = 4576; cin = 0;
#10 a = 39782; b = 6057; cin = 1;
#10 a = 43191; b = 64241; cin = 0;
#10 a = 62418; b = 2553; cin = 1;
#10 a = 53337; b = 22302; cin = 1;
#10 a = 34210; b = 9078; cin = 1;
#10 a = 56791; b = 48407; cin = 0;
#10 a = 34797; b = 24800; cin = 1;
#10 a = 21071; b = 16921; cin = 1;
#10 a = 26346; b = 66154; cin = 0;
#10 a = 18089; b = 35275; cin = 0;
#10 a = 31341; b = 51409; cin = 1;
#10 a = 10074; b = 24600; cin = 0;
#10 a = 1197; b = 63371; cin = 1;
#10 a = 33722; b = 46708; cin = 1;
#10 a = 48403; b = 57270; cin = 0;
#10 a = 33683; b = 44061; cin = 1;
#10 a = 57579; b = 55210; cin = 1;
#10 a = 5702; b = 6282; cin = 0;
#10 a = 50537; b = 32628; cin = 0;
#10 a = 22455; b = 27069; cin = 1;
#10 a = 45301; b = 34763; cin = 0;
#10 a = 50556; b = 44837; cin = 1;
#10 a = 50052; b = 22386; cin = 0;
#10 a = 28453; b = 32461; cin = 0;
#10 a = 29156; b = 10864; cin = 1;
#10 a = 38938; b = 44547; cin = 0;
#10 a = 3479; b = 32126; cin = 1;
#10 a = 39173; b = 14180; cin = 1;
#10 a = 21787; b = 41069; cin = 1;
#10 a = 46908; b = 39876; cin = 1;
#10 a = 13655; b = 15177; cin = 0;
#10 a = 8164; b = 42085; cin = 1;
#10 a = 3625; b = 68489; cin = 0;
#10 a = 38809; b = 26942; cin = 1;
#10 a = 50701; b = 56099; cin = 1;
#10 a = 49864; b = 1389; cin = 1;
#10 a = 69441; b = 51221; cin = 1;
#10 a = 4228; b = 20394; cin = 0;
#10 a = 15297; b = 18533; cin = 1;
#10 a = 11698; b = 65441; cin = 0;
#10 a = 35169; b = 55449; cin = 1;
#10 a = 69755; b = 39965; cin = 1;
#10 a = 55531; b = 19942; cin = 0;
#10 a = 63693; b = 58751; cin = 1;
#10 a = 10668; b = 39452; cin = 0;
#10 a = 62155; b = 65669; cin = 1;
#10 a = 64542; b = 65110; cin = 0;
#10 a = 5408; b = 69338; cin = 0;
#10 a = 30454; b = 60987; cin = 0;
#10 a = 2921; b = 2685; cin = 1;
#10 a = 15265; b = 37855; cin = 0;
#10 a = 19139; b = 13962; cin = 1;
#10 a = 41450; b = 69493; cin = 1;
#10 a = 15898; b = 63186; cin = 0;
#10 a = 63641; b = 50206; cin = 1;
#10 a = 3835; b = 42362; cin = 0;
#10 a = 15419; b = 13256; cin = 0;
#10 a = 8223; b = 18664; cin = 0;
#10 a = 67774; b = 49118; cin = 1;
#10 a = 5858; b = 28392; cin = 0;
#10 a = 9383; b = 43657; cin = 1;
#10 a = 21062; b = 39148; cin = 0;
#10 a = 2705; b = 10598; cin = 1;
#10 a = 50643; b = 2849; cin = 0;
#10 a = 17331; b = 66490; cin = 0;
#10 a = 69824; b = 46678; cin = 0;
#10 a = 47986; b = 62097; cin = 1;
#10 a = 21258; b = 320; cin = 1;
#10 a = 16572; b = 68094; cin = 0;
#10 a = 26521; b = 3952; cin = 0;
#10 a = 15508; b = 59688; cin = 1;
#10 a = 18701; b = 10750; cin = 0;
#10 a = 35857; b = 59807; cin = 0;
#10 a = 28859; b = 40450; cin = 1;
#10 a = 15047; b = 57782; cin = 0;
#10 a = 51441; b = 33958; cin = 0;
#10 a = 12902; b = 11945; cin = 1;
#10 a = 11267; b = 9555; cin = 1;
#10 a = 4648; b = 26128; cin = 0;
#10 a = 23500; b = 29001; cin = 0;
#10 a = 744; b = 20861; cin = 0;
#10 a = 67998; b = 39563; cin = 0;
#10 a = 10752; b = 51772; cin = 0;
#10 a = 57752; b = 10631; cin = 0;
#10 a = 13954; b = 25678; cin = 0;
#10 a = 12998; b = 53472; cin = 1;
#10 a = 12368; b = 66374; cin = 0;
#10 a = 50187; b = 53993; cin = 1;
#10 a = 64678; b = 58641; cin = 1;
#10 a = 7264; b = 58494; cin = 1;
#10 a = 155; b = 35590; cin = 0;
#10 a = 29085; b = 33588; cin = 1;
#10 a = 45118; b = 20692; cin = 0;
#10 a = 50958; b = 8445; cin = 1;
#10 a = 27248; b = 68751; cin = 0;
#10 a = 14025; b = 11749; cin = 0;
#10 a = 58408; b = 469; cin = 0;
#10 a = 21088; b = 27008; cin = 1;
#10 a = 16027; b = 21686; cin = 0;
#10 a = 60743; b = 5303; cin = 0;
#10 a = 17164; b = 51810; cin = 1;
#10 a = 18094; b = 57247; cin = 1;
#10 a = 34940; b = 32365; cin = 0;
#10 a = 9910; b = 13323; cin = 1;
#10 a = 65511; b = 16924; cin = 0;
#10 a = 6791; b = 30949; cin = 1;
#10 a = 24247; b = 65709; cin = 0;
#10 a = 61725; b = 63149; cin = 0;
#10 a = 59548; b = 9176; cin = 0;
#10 a = 22365; b = 69919; cin = 1;
#10 a = 43675; b = 63435; cin = 1;
#10 a = 30576; b = 57882; cin = 1;
#10 a = 3770; b = 22822; cin = 0;
#10 a = 21304; b = 9084; cin = 0;
#10 a = 69987; b = 4595; cin = 0;
#10 a = 47421; b = 57739; cin = 1;
#10 a = 12956; b = 11986; cin = 0;
#10 a = 48960; b = 50064; cin = 1;
#10 a = 18324; b = 15964; cin = 1;
#10 a = 32078; b = 38329; cin = 1;
#10 a = 4784; b = 58357; cin = 0;
#10 a = 52003; b = 65285; cin = 0;
#10 a = 16470; b = 69055; cin = 0;
#10 a = 13303; b = 66711; cin = 0;
#10 a = 69811; b = 66698; cin = 0;
#10 a = 3243; b = 44119; cin = 1;
#10 a = 13976; b = 57075; cin = 1;
#10 a = 20418; b = 12387; cin = 1;
#10 a = 43657; b = 7063; cin = 0;
#10 a = 52424; b = 39142; cin = 1;
#10 a = 37463; b = 20278; cin = 0;
#10 a = 15938; b = 48633; cin = 0;
#10 a = 52294; b = 65104; cin = 1;
#10 a = 17825; b = 8407; cin = 1;
#10 a = 62439; b = 8218; cin = 1;
#10 a = 18001; b = 57813; cin = 1;
#10 a = 7654; b = 1789; cin = 0;
#10 a = 55646; b = 68559; cin = 0;
#10 a = 13701; b = 42216; cin = 1;
#10 a = 34073; b = 992; cin = 1;
#10 a = 22775; b = 38456; cin = 1;
#10 a = 46185; b = 30746; cin = 1;
#10 a = 41233; b = 13040; cin = 1;
#10 a = 35337; b = 30865; cin = 0;
#10 a = 26152; b = 69657; cin = 0;
#10 a = 60017; b = 64010; cin = 1;
#10 a = 44354; b = 1665; cin = 0;
#10 a = 15767; b = 33663; cin = 1;
#10 a = 45919; b = 47364; cin = 1;
#10 a = 13134; b = 11438; cin = 1;
#10 a = 65844; b = 10565; cin = 1;
#10 a = 68831; b = 33102; cin = 1;
#10 a = 50452; b = 4336; cin = 0;
#10 a = 3529; b = 39673; cin = 1;
#10 a = 35013; b = 42177; cin = 0;
#10 a = 51067; b = 32194; cin = 1;
#10 a = 54934; b = 6549; cin = 0;
#10 a = 13294; b = 68668; cin = 1;
#10 a = 40213; b = 44587; cin = 1;
#10 a = 39348; b = 34073; cin = 1;
#10 a = 15828; b = 29917; cin = 0;
#10 a = 30763; b = 5101; cin = 1;
#10 a = 52797; b = 31905; cin = 1;
#10 a = 17871; b = 35435; cin = 0;
#10 a = 60162; b = 448; cin = 1;
#10 a = 32111; b = 27868; cin = 1;
#10 a = 68070; b = 59154; cin = 0;
#10 a = 12046; b = 2449; cin = 0;
#10 a = 59685; b = 42662; cin = 1;
#10 a = 61040; b = 58363; cin = 1;
#10 a = 50186; b = 4191; cin = 0;
#10 a = 49896; b = 11306; cin = 1;
#10 a = 12709; b = 40455; cin = 1;
#10 a = 49858; b = 58326; cin = 0;
#10 a = 56680; b = 48489; cin = 0;
#10 a = 12031; b = 56952; cin = 0;
#10 a = 69577; b = 55022; cin = 1;
#10 a = 40023; b = 43420; cin = 0;
#10 a = 55490; b = 9457; cin = 0;
#10 a = 45543; b = 46849; cin = 1;
#10 a = 22374; b = 27035; cin = 0;
#10 a = 52771; b = 6932; cin = 1;
#10 a = 64620; b = 19641; cin = 0;
#10 a = 38375; b = 69500; cin = 1;
#10 a = 47565; b = 32532; cin = 0;
#10 a = 33556; b = 44564; cin = 0;
#10 a = 47414; b = 44141; cin = 0;
#10 a = 50427; b = 14164; cin = 0;
#10 a = 32241; b = 46006; cin = 1;
#10 a = 33070; b = 67902; cin = 0;
#10 a = 22261; b = 20276; cin = 0;
#10 a = 61996; b = 3047; cin = 0;
#10 a = 43037; b = 44020; cin = 1;
#10 a = 40885; b = 58747; cin = 1;
#10 a = 3412; b = 36313; cin = 0;
#10 a = 14428; b = 46221; cin = 0;
#10 a = 58748; b = 23635; cin = 1;
#10 a = 64442; b = 50415; cin = 1;
#10 a = 43556; b = 59008; cin = 0;
#10 a = 8479; b = 22078; cin = 0;
#10 a = 20252; b = 44340; cin = 0;
#10 a = 59060; b = 36336; cin = 0;
#10 a = 34800; b = 9373; cin = 0;
#10 a = 30181; b = 26610; cin = 1;
#10 a = 1415; b = 30023; cin = 0;
#10 a = 5181; b = 20803; cin = 1;
#10 a = 53511; b = 9552; cin = 1;
#10 a = 52334; b = 50346; cin = 0;
#10 a = 41673; b = 255; cin = 0;
#10 a = 30667; b = 8734; cin = 1;
#10 a = 63915; b = 28986; cin = 1;
#10 a = 23792; b = 64398; cin = 1;
#10 a = 56716; b = 29198; cin = 0;
#10 a = 40012; b = 35732; cin = 0;
#10 a = 35703; b = 37147; cin = 1;
#10 a = 20412; b = 18680; cin = 1;
#10 a = 51341; b = 48543; cin = 1;
#10 a = 35906; b = 7229; cin = 1;
#10 a = 47238; b = 48902; cin = 0;
#10 a = 23931; b = 55922; cin = 1;
#10 a = 46350; b = 26189; cin = 1;
#10 a = 19461; b = 49981; cin = 0;
#10 a = 28908; b = 36697; cin = 0;
#10 a = 24080; b = 6709; cin = 0;
#10 a = 22214; b = 18765; cin = 1;
#10 a = 50372; b = 15529; cin = 1;
#10 a = 5685; b = 66870; cin = 0;
#10 a = 40550; b = 32777; cin = 1;
#10 a = 32113; b = 56367; cin = 0;
#10 a = 23932; b = 10298; cin = 0;
#10 a = 837; b = 33000; cin = 1;
#10 a = 53080; b = 52461; cin = 1;
#10 a = 53370; b = 57721; cin = 0;
#10 a = 59211; b = 58153; cin = 0;
#10 a = 30783; b = 10368; cin = 1;
#10 a = 15855; b = 37092; cin = 0;
#10 a = 65958; b = 19129; cin = 0;
#10 a = 957; b = 36031; cin = 1;
#10 a = 13184; b = 68144; cin = 1;
#10 a = 4314; b = 68428; cin = 1;
#10 a = 51366; b = 45617; cin = 0;
#10 a = 54608; b = 28698; cin = 1;
#10 a = 14183; b = 12068; cin = 1;
#10 a = 10455; b = 47631; cin = 0;
#10 a = 59789; b = 54767; cin = 0;
#10 a = 57888; b = 622; cin = 0;
#10 a = 47868; b = 42932; cin = 1;
#10 a = 58367; b = 43889; cin = 0;
#10 a = 54346; b = 57074; cin = 1;
#10 a = 36693; b = 37740; cin = 1;
#10 a = 29339; b = 19107; cin = 1;
#10 a = 31337; b = 50067; cin = 1;
#10 a = 15796; b = 40602; cin = 1;
#10 a = 57977; b = 51057; cin = 1;
#10 a = 64664; b = 17199; cin = 0;
#10 a = 11718; b = 5087; cin = 0;
#10 a = 42217; b = 29308; cin = 0;
#10 a = 21844; b = 64027; cin = 0;
#10 a = 37503; b = 48373; cin = 0;
#10 a = 27658; b = 15067; cin = 0;
#10 a = 62593; b = 44406; cin = 1;
#10 a = 3146; b = 52095; cin = 0;
#10 a = 18749; b = 44243; cin = 0;
#10 a = 46421; b = 32221; cin = 0;
#10 a = 28076; b = 3237; cin = 1;
#10 a = 18146; b = 14955; cin = 0;
#10 a = 31542; b = 33524; cin = 0;
#10 a = 64222; b = 55369; cin = 1;
#10 a = 792; b = 69224; cin = 1;
#10 a = 40788; b = 26882; cin = 0;
#10 a = 24877; b = 65827; cin = 0;
#10 a = 28072; b = 45326; cin = 1;
#10 a = 11335; b = 64075; cin = 0;
#10 a = 11551; b = 40496; cin = 1;
#10 a = 62825; b = 68572; cin = 0;
#10 a = 61298; b = 63070; cin = 0;
#10 a = 17563; b = 964; cin = 0;
#10 a = 26783; b = 65187; cin = 1;
#10 a = 6383; b = 65979; cin = 1;
#10 a = 34356; b = 13120; cin = 1;
#10 a = 7396; b = 37997; cin = 1;
#10 a = 24842; b = 66069; cin = 1;
#10 a = 47087; b = 7404; cin = 0;
#10 a = 67223; b = 65308; cin = 1;
#10 a = 2285; b = 58133; cin = 1;
#10 a = 34231; b = 25784; cin = 0;
#10 a = 33837; b = 43347; cin = 0;
#10 a = 20616; b = 46482; cin = 1;
#10 a = 39115; b = 52865; cin = 1;
#10 a = 56839; b = 17221; cin = 1;
#10 a = 7796; b = 24617; cin = 0;
#10 a = 24581; b = 25811; cin = 1;
#10 a = 63044; b = 49250; cin = 0;
#10 a = 25583; b = 46474; cin = 0;
#10 a = 4970; b = 25111; cin = 1;
#10 a = 52929; b = 59342; cin = 1;
#10 a = 311; b = 23180; cin = 0;
#10 a = 18658; b = 20148; cin = 1;
#10 a = 32191; b = 59263; cin = 0;
#10 a = 18056; b = 22454; cin = 0;
#10 a = 17041; b = 30251; cin = 1;
#10 a = 54023; b = 31184; cin = 1;
#10 a = 63427; b = 24229; cin = 1;
#10 a = 10235; b = 26164; cin = 1;
#10 a = 68703; b = 31134; cin = 0;
#10 a = 21656; b = 14063; cin = 1;
#10 a = 394; b = 60727; cin = 1;
#10 a = 22478; b = 9385; cin = 1;
#10 a = 67397; b = 41576; cin = 0;
#10 a = 1534; b = 35985; cin = 1;
#10 a = 69244; b = 53026; cin = 0;
#10 a = 67923; b = 13402; cin = 0;
#10 a = 22414; b = 6829; cin = 1;
#10 a = 26156; b = 63416; cin = 1;
#10 a = 29075; b = 38471; cin = 1;
#10 a = 10754; b = 60127; cin = 1;
#10 a = 28127; b = 60521; cin = 0;
#10 a = 45032; b = 59352; cin = 1;
#10 a = 12085; b = 33101; cin = 1;
#10 a = 14753; b = 10987; cin = 0;
#10 a = 39876; b = 10231; cin = 1;
#10 a = 1602; b = 54507; cin = 1;
#10 a = 64513; b = 6921; cin = 0;
#10 a = 58004; b = 9429; cin = 0;
#10 a = 7660; b = 38505; cin = 1;
#10 a = 34801; b = 25611; cin = 0;
#10 a = 52358; b = 30090; cin = 0;
#10 a = 60642; b = 51474; cin = 0;
#10 a = 54663; b = 39911; cin = 1;
#10 a = 20261; b = 31016; cin = 1;
#10 a = 21843; b = 893; cin = 0;
#10 a = 52804; b = 48847; cin = 1;
#10 a = 27167; b = 43360; cin = 1;
#10 a = 8359; b = 7717; cin = 0;
#10 a = 52967; b = 61729; cin = 1;
#10 a = 42398; b = 2882; cin = 0;
#10 a = 21957; b = 55241; cin = 0;
#10 a = 62037; b = 22235; cin = 0;
#10 a = 67821; b = 53251; cin = 1;
#10 a = 60354; b = 3512; cin = 0;
#10 a = 40227; b = 1707; cin = 1;
#10 a = 6684; b = 30864; cin = 0;
#10 a = 27647; b = 58031; cin = 1;
#10 a = 55532; b = 42743; cin = 0;
#10 a = 69199; b = 2062; cin = 1;
#10 a = 27722; b = 20813; cin = 1;
#10 a = 11857; b = 42770; cin = 0;
#10 a = 2433; b = 11159; cin = 0;
#10 a = 20836; b = 8980; cin = 1;
#10 a = 9149; b = 45686; cin = 1;
#10 a = 28479; b = 62266; cin = 0;
#10 a = 1406; b = 45302; cin = 0;
#10 a = 46829; b = 2949; cin = 0;
#10 a = 41964; b = 34834; cin = 1;
#10 a = 44816; b = 10385; cin = 1;
#10 a = 39397; b = 38107; cin = 0;
#10 a = 13212; b = 26316; cin = 0;
#10 a = 42269; b = 5102; cin = 1;
#10 a = 69913; b = 25938; cin = 1;
#10 a = 10808; b = 11439; cin = 0;
#10 a = 47919; b = 39919; cin = 0;
#10 a = 16737; b = 41325; cin = 0;
#10 a = 62772; b = 64506; cin = 1;
#10 a = 26838; b = 36470; cin = 1;
#10 a = 56351; b = 57638; cin = 0;
#10 a = 41574; b = 3387; cin = 0;
#10 a = 23963; b = 16600; cin = 0;
#10 a = 49121; b = 58869; cin = 0;
#10 a = 15439; b = 35134; cin = 0;
#10 a = 37088; b = 22294; cin = 0;
#10 a = 58072; b = 213; cin = 1;
#10 a = 47674; b = 16950; cin = 0;
#10 a = 12578; b = 9722; cin = 1;
#10 a = 26784; b = 12912; cin = 1;
#10 a = 5823; b = 45615; cin = 0;
#10 a = 41600; b = 63542; cin = 1;
#10 a = 21836; b = 17505; cin = 1;
#10 a = 28388; b = 42978; cin = 0;
#10 a = 16395; b = 34769; cin = 0;
#10 a = 6691; b = 1858; cin = 0;
#10 a = 8427; b = 59930; cin = 1;
#10 a = 26434; b = 13957; cin = 0;
#10 a = 62119; b = 2887; cin = 0;
#10 a = 68662; b = 29671; cin = 1;
#10 a = 41675; b = 35495; cin = 0;
#10 a = 25031; b = 53447; cin = 0;
#10 a = 35423; b = 5283; cin = 1;
#10 a = 38766; b = 10023; cin = 0;
#10 a = 7331; b = 26418; cin = 1;
#10 a = 57381; b = 9462; cin = 1;
#10 a = 13374; b = 64241; cin = 0;
#10 a = 15931; b = 67028; cin = 1;
#10 a = 11791; b = 59147; cin = 0;
#10 a = 17374; b = 34161; cin = 0;
#10 a = 58573; b = 52188; cin = 1;
#10 a = 5387; b = 7220; cin = 0;
#10 a = 39392; b = 42643; cin = 1;
#10 a = 43605; b = 57761; cin = 0;
#10 a = 44445; b = 41444; cin = 1;
#10 a = 56407; b = 28826; cin = 1;
#10 a = 226; b = 18552; cin = 0;
#10 a = 50328; b = 10835; cin = 0;
#10 a = 44387; b = 22627; cin = 1;
#10 a = 41334; b = 16353; cin = 0;
#10 a = 44304; b = 4926; cin = 1;
#10 a = 12769; b = 56665; cin = 1;
#10 a = 11033; b = 26057; cin = 0;
#10 a = 14580; b = 46015; cin = 1;
#10 a = 28150; b = 66812; cin = 0;
#10 a = 44491; b = 53219; cin = 0;
#10 a = 46646; b = 29798; cin = 0;
#10 a = 43043; b = 10126; cin = 1;
#10 a = 36467; b = 30866; cin = 0;
#10 a = 19039; b = 48552; cin = 1;
#10 a = 12123; b = 22856; cin = 1;
#10 a = 57396; b = 11977; cin = 1;
#10 a = 16241; b = 69362; cin = 0;
#10 a = 41377; b = 13942; cin = 1;
#10 a = 6979; b = 18444; cin = 0;
#10 a = 14025; b = 62936; cin = 1;
#10 a = 26249; b = 39582; cin = 1;
#10 a = 57025; b = 58977; cin = 0;
#10 a = 51340; b = 25445; cin = 0;
#10 a = 68283; b = 20836; cin = 0;
#10 a = 7930; b = 9311; cin = 0;
#10 a = 68856; b = 43060; cin = 1;
#10 a = 46447; b = 59301; cin = 1;
#10 a = 50095; b = 30679; cin = 1;
#10 a = 6111; b = 14010; cin = 1;
#10 a = 28939; b = 28035; cin = 1;
#10 a = 11338; b = 54284; cin = 0;
#10 a = 23536; b = 17661; cin = 1;
#10 a = 45860; b = 69001; cin = 0;
#10 a = 5402; b = 67284; cin = 0;
#10 a = 13496; b = 51567; cin = 0;
#10 a = 20798; b = 50423; cin = 0;
#10 a = 16429; b = 26870; cin = 1;
#10 a = 35070; b = 53317; cin = 0;
#10 a = 44005; b = 59428; cin = 0;
#10 a = 1384; b = 64719; cin = 1;
#10 a = 68052; b = 6058; cin = 1;
#10 a = 10654; b = 5946; cin = 0;
#10 a = 35881; b = 28158; cin = 0;
#10 a = 62906; b = 33560; cin = 0;
#10 a = 40766; b = 23408; cin = 1;
#10 a = 4290; b = 20558; cin = 0;
#10 a = 34522; b = 36987; cin = 0;
#10 a = 54056; b = 48409; cin = 0;
#10 a = 10620; b = 68766; cin = 0;
#10 a = 51195; b = 150; cin = 0;
#10 a = 49804; b = 44554; cin = 0;
#10 a = 9050; b = 55208; cin = 0;
#10 a = 55956; b = 67442; cin = 0;
#10 a = 31864; b = 36700; cin = 0;
#10 a = 5057; b = 53818; cin = 0;
#10 a = 6168; b = 58109; cin = 0;
#10 a = 34055; b = 22631; cin = 1;
#10 a = 42459; b = 6687; cin = 0;
#10 a = 10533; b = 63660; cin = 0;
#10 a = 14388; b = 44855; cin = 0;
#10 a = 59314; b = 1011; cin = 1;
#10 a = 16650; b = 10061; cin = 1;
#10 a = 49932; b = 66018; cin = 1;
#10 a = 41372; b = 4234; cin = 1;
#10 a = 66372; b = 9291; cin = 0;
#10 a = 67484; b = 61812; cin = 1;
#10 a = 19154; b = 25867; cin = 0;
#10 a = 54163; b = 44678; cin = 0;
#10 a = 21229; b = 31564; cin = 0;
#10 a = 33413; b = 22304; cin = 1;
#10 a = 22099; b = 57970; cin = 0;
#10 a = 31692; b = 4620; cin = 0;
#10 a = 26494; b = 54552; cin = 0;
#10 a = 65089; b = 25924; cin = 0;
#10 a = 385; b = 68648; cin = 0;
#10 a = 59499; b = 66132; cin = 0;
#10 a = 36722; b = 61638; cin = 1;
#10 a = 12928; b = 45801; cin = 1;
#10 a = 42174; b = 43382; cin = 1;
#10 a = 65080; b = 53147; cin = 1;
#10 a = 39193; b = 51598; cin = 1;
#10 a = 14318; b = 13291; cin = 1;
#10 a = 45856; b = 16137; cin = 1;
#10 a = 49764; b = 11226; cin = 1;
#10 a = 34258; b = 11611; cin = 1;
#10 a = 28044; b = 1110; cin = 1;
#10 a = 59994; b = 14184; cin = 1;
#10 a = 24163; b = 3465; cin = 0;
#10 a = 33011; b = 45639; cin = 0;
#10 a = 49774; b = 17072; cin = 1;
#10 a = 65194; b = 56265; cin = 0;
#10 a = 68583; b = 583; cin = 1;
#10 a = 6593; b = 22791; cin = 0;
#10 a = 45506; b = 48907; cin = 0;
#10 a = 40344; b = 13166; cin = 0;
#10 a = 33829; b = 17562; cin = 0;
#10 a = 46151; b = 7557; cin = 1;
#10 a = 50110; b = 31720; cin = 0;
#10 a = 29871; b = 64731; cin = 1;
#10 a = 5717; b = 20858; cin = 1;
#10 a = 34711; b = 62404; cin = 1;
#10 a = 45303; b = 60987; cin = 0;
#10 a = 45538; b = 43932; cin = 0;
#10 a = 61910; b = 19439; cin = 1;
#10 a = 19508; b = 36135; cin = 1;
#10 a = 58718; b = 46316; cin = 0;
#10 a = 5391; b = 22467; cin = 1;
#10 a = 36248; b = 2578; cin = 1;
#10 a = 570; b = 8801; cin = 1;
#10 a = 56883; b = 14518; cin = 1;
#10 a = 36621; b = 49229; cin = 1;
#10 a = 26272; b = 884; cin = 0;
#10 a = 62858; b = 46422; cin = 1;
#10 a = 28588; b = 38332; cin = 0;
#10 a = 43226; b = 57841; cin = 1;
#10 a = 1029; b = 46559; cin = 1;
#10 a = 22747; b = 51950; cin = 1;
#10 a = 52022; b = 18198; cin = 1;
#10 a = 43018; b = 65120; cin = 0;
#10 a = 5097; b = 28356; cin = 0;
#10 a = 34386; b = 64977; cin = 0;
#10 a = 32431; b = 21249; cin = 0;
#10 a = 21463; b = 60459; cin = 1;
#10 a = 54428; b = 65400; cin = 1;
#10 a = 59536; b = 38626; cin = 0;
#10 a = 30779; b = 16007; cin = 0;
#10 a = 1987; b = 15107; cin = 0;
#10 a = 18366; b = 67129; cin = 1;
#10 a = 37323; b = 16499; cin = 1;
#10 a = 41433; b = 21596; cin = 1;
#10 a = 36413; b = 32334; cin = 0;
#10 a = 56975; b = 64765; cin = 1;
#10 a = 8422; b = 62581; cin = 1;
#10 a = 6291; b = 23361; cin = 1;
#10 a = 18844; b = 12898; cin = 1;
#10 a = 19239; b = 43677; cin = 0;
#10 a = 42545; b = 22016; cin = 1;
#10 a = 24153; b = 40382; cin = 1;
#10 a = 23960; b = 54057; cin = 0;
#10 a = 65240; b = 1842; cin = 1;
#10 a = 64875; b = 38256; cin = 1;
#10 a = 35840; b = 1583; cin = 1;
#10 a = 4405; b = 10005; cin = 0;
#10 a = 33430; b = 62648; cin = 1;
#10 a = 34207; b = 11493; cin = 1;
#10 a = 3610; b = 7084; cin = 1;
#10 a = 35373; b = 25981; cin = 1;
#10 a = 12242; b = 50134; cin = 0;
#10 a = 56241; b = 50447; cin = 1;
#10 a = 23092; b = 45687; cin = 0;
#10 a = 11539; b = 16914; cin = 0;
#10 a = 8672; b = 29106; cin = 1;
#10 a = 46923; b = 33512; cin = 1;
#10 a = 7755; b = 43294; cin = 1;
#10 a = 61949; b = 7502; cin = 0;
#10 a = 35392; b = 57464; cin = 0;
#10 a = 52513; b = 22837; cin = 1;
#10 a = 21651; b = 11432; cin = 0;
#10 a = 7523; b = 44025; cin = 1;
#10 a = 23804; b = 67117; cin = 0;
#10 a = 65576; b = 55008; cin = 0;
#10 a = 28308; b = 63681; cin = 1;
#10 a = 16272; b = 16956; cin = 1;
#10 a = 60593; b = 24712; cin = 1;
#10 a = 27562; b = 63013; cin = 1;
#10 a = 52377; b = 28405; cin = 0;
#10 a = 60627; b = 57271; cin = 1;
#10 a = 24859; b = 8922; cin = 1;
#10 a = 39225; b = 62797; cin = 1;
#10 a = 10390; b = 16601; cin = 0;
#10 a = 27242; b = 58530; cin = 1;
#10 a = 13712; b = 16838; cin = 0;
#10 a = 52937; b = 33110; cin = 0;
#10 a = 32026; b = 55; cin = 0;
#10 a = 30762; b = 3970; cin = 1;
#10 a = 36999; b = 56347; cin = 1;
#10 a = 7053; b = 23326; cin = 0;
#10 a = 69945; b = 48185; cin = 0;
#10 a = 50620; b = 63762; cin = 1;
#10 a = 5321; b = 4152; cin = 0;
#10 a = 27140; b = 7746; cin = 0;
#10 a = 10319; b = 21459; cin = 1;
#10 a = 33531; b = 50748; cin = 1;
#10 a = 27347; b = 59127; cin = 1;
#10 a = 68580; b = 19889; cin = 1;
#10 a = 56473; b = 33240; cin = 0;
#10 a = 25476; b = 40294; cin = 0;
#10 a = 51750; b = 40239; cin = 0;
#10 a = 16946; b = 20859; cin = 0;
#10 a = 21291; b = 2533; cin = 1;
#10 a = 42238; b = 6025; cin = 1;
#10 a = 28066; b = 16344; cin = 0;
#10 a = 30733; b = 26227; cin = 1;
#10 a = 19215; b = 53574; cin = 0;
#10 a = 31400; b = 28506; cin = 1;
#10 a = 23907; b = 14980; cin = 1;
#10 a = 2761; b = 16808; cin = 1;
#10 a = 51293; b = 68559; cin = 0;
#10 a = 8011; b = 15505; cin = 0;
#10 a = 52140; b = 13149; cin = 1;
#10 a = 53125; b = 55387; cin = 0;
#10 a = 15504; b = 59805; cin = 0;
#10 a = 22047; b = 66891; cin = 1;
#10 a = 32986; b = 16106; cin = 1;
#10 a = 55756; b = 23858; cin = 0;
#10 a = 52063; b = 47765; cin = 0;
#10 a = 34314; b = 26878; cin = 0;
#10 a = 56860; b = 8171; cin = 1;
#10 a = 49644; b = 62535; cin = 1;
#10 a = 39640; b = 21027; cin = 0;
#10 a = 8521; b = 4152; cin = 1;
#10 a = 7075; b = 66008; cin = 0;
#10 a = 44677; b = 18055; cin = 1;
#10 a = 62154; b = 27393; cin = 1;
#10 a = 15910; b = 13149; cin = 1;
#10 a = 21820; b = 41564; cin = 0;
#10 a = 19062; b = 5879; cin = 0;
#10 a = 9464; b = 62739; cin = 0;
#10 a = 22074; b = 18735; cin = 1;
#10 a = 26541; b = 34728; cin = 0;
#10 a = 20509; b = 43249; cin = 0;
#10 a = 69864; b = 26677; cin = 0;
#10 a = 39024; b = 1354; cin = 0;
#10 a = 51428; b = 39861; cin = 1;
#10 a = 56289; b = 55771; cin = 1;
#10 a = 15009; b = 53943; cin = 1;
#10 a = 21493; b = 49357; cin = 0;
#10 a = 7560; b = 58821; cin = 1;
#10 a = 1798; b = 10895; cin = 1;
#10 a = 58571; b = 13788; cin = 1;
#10 a = 66371; b = 34297; cin = 0;
#10 a = 8323; b = 34161; cin = 1;
#10 a = 62635; b = 49538; cin = 0;
#10 a = 65003; b = 7318; cin = 1;
#10 a = 1117; b = 39959; cin = 0;
#10 a = 44028; b = 54968; cin = 1;
#10 a = 11207; b = 52814; cin = 0;
#10 a = 54266; b = 60374; cin = 1;
#10 a = 66415; b = 62172; cin = 1;
#10 a = 50948; b = 50743; cin = 1;
#10 a = 22913; b = 47114; cin = 1;
#10 a = 38128; b = 31789; cin = 0;
#10 a = 10019; b = 776; cin = 0;
#10 a = 5969; b = 65780; cin = 0;
#10 a = 41780; b = 66897; cin = 0;
#10 a = 39714; b = 17277; cin = 0;
#10 a = 21591; b = 28484; cin = 0;
#10 a = 29177; b = 59102; cin = 0;
#10 a = 49233; b = 55518; cin = 0;
#10 a = 32888; b = 12818; cin = 1;
#10 a = 30331; b = 35732; cin = 1;
#10 a = 38424; b = 3860; cin = 0;
#10 a = 57031; b = 60231; cin = 1;
#10 a = 31527; b = 66201; cin = 1;
#10 a = 13342; b = 37981; cin = 0;
#10 a = 35116; b = 54048; cin = 1;
#10 a = 18210; b = 51991; cin = 1;
#10 a = 54119; b = 11169; cin = 0;
#10 a = 10401; b = 36754; cin = 0;
#10 a = 5208; b = 69642; cin = 0;
#10 a = 27109; b = 6325; cin = 0;
#10 a = 26125; b = 21102; cin = 0;
#10 a = 9633; b = 8133; cin = 0;
#10 a = 17566; b = 16012; cin = 1;
#10 a = 67631; b = 29354; cin = 0;
#10 a = 20945; b = 64470; cin = 0;
#10 a = 61536; b = 59033; cin = 0;
#10 a = 13316; b = 43152; cin = 1;
#10 a = 24198; b = 29905; cin = 1;
#10 a = 20598; b = 11465; cin = 1;
#10 a = 29816; b = 14927; cin = 0;
#10 a = 51119; b = 17404; cin = 0;
#10 a = 6281; b = 27037; cin = 1;
#10 a = 68027; b = 20956; cin = 0;
#10 a = 55974; b = 18587; cin = 0;
#10 a = 58255; b = 15885; cin = 1;
#10 a = 44583; b = 53773; cin = 0;
#10 a = 59255; b = 67089; cin = 0;
#10 a = 15096; b = 21287; cin = 1;
#10 a = 54043; b = 41885; cin = 1;
#10 a = 68984; b = 48054; cin = 0;
#10 a = 20251; b = 29173; cin = 0;
#10 a = 38971; b = 11806; cin = 1;
#10 a = 42177; b = 9834; cin = 1;
#10 a = 15043; b = 65808; cin = 1;
#10 a = 63615; b = 54063; cin = 0;
#10 a = 13010; b = 4999; cin = 1;
#10 a = 67790; b = 40606; cin = 1;
#10 a = 49370; b = 32055; cin = 0;
#10 a = 13560; b = 16098; cin = 0;
#10 a = 59215; b = 61435; cin = 0;
#10 a = 49797; b = 11686; cin = 1;
#10 a = 34135; b = 27009; cin = 1;
#10 a = 69158; b = 69186; cin = 1;
#10 a = 31490; b = 60581; cin = 0;
#10 a = 12409; b = 30549; cin = 1;
#10 a = 55565; b = 19911; cin = 0;
#10 a = 58846; b = 17702; cin = 1;
#10 a = 59217; b = 43424; cin = 0;
#10 a = 57228; b = 56984; cin = 0;
#10 a = 3476; b = 22551; cin = 1;
#10 a = 44130; b = 48700; cin = 1;
#10 a = 43957; b = 12835; cin = 1;
#10 a = 55590; b = 11994; cin = 1;
#10 a = 53410; b = 43484; cin = 1;
#10 a = 47038; b = 32245; cin = 0;
#10 a = 24729; b = 64162; cin = 1;
#10 a = 30124; b = 53008; cin = 1;
#10 a = 6125; b = 42226; cin = 0;
#10 a = 60533; b = 5806; cin = 0;
#10 a = 61039; b = 55634; cin = 0;
#10 a = 29333; b = 6116; cin = 0;
#10 a = 9312; b = 50073; cin = 0;
#10 a = 62653; b = 12015; cin = 0;
#10 a = 21533; b = 65425; cin = 0;
#10 a = 40994; b = 42463; cin = 1;
#10 a = 21004; b = 43545; cin = 1;
#10 a = 67277; b = 50021; cin = 1;
#10 a = 37605; b = 32498; cin = 1;
#10 a = 5005; b = 23031; cin = 1;
#10 a = 5741; b = 14070; cin = 1;
#10 a = 5381; b = 43403; cin = 1;
#10 a = 53722; b = 29068; cin = 0;
#10 a = 44898; b = 68073; cin = 0;
#10 a = 48068; b = 19606; cin = 1;
#10 a = 47426; b = 60600; cin = 1;
#10 a = 9029; b = 57956; cin = 0;
#10 a = 34794; b = 31586; cin = 1;
#10 a = 19919; b = 69191; cin = 1;
#10 a = 47271; b = 50548; cin = 0;
#10 a = 56780; b = 32641; cin = 0;
#10 a = 51924; b = 38023; cin = 0;
#10 a = 29535; b = 21745; cin = 0;
#10 a = 57220; b = 66643; cin = 1;
#10 a = 26920; b = 21063; cin = 0;
#10 a = 14749; b = 68489; cin = 0;
#10 a = 21394; b = 53870; cin = 1;
#10 a = 1584; b = 18664; cin = 1;
#10 a = 8147; b = 14935; cin = 0;
#10 a = 23560; b = 62206; cin = 0;
#10 a = 15652; b = 25339; cin = 1;
#10 a = 44519; b = 7263; cin = 0;
#10 a = 23141; b = 36798; cin = 1;
#10 a = 30831; b = 24018; cin = 0;
#10 a = 36594; b = 27290; cin = 1;
#10 a = 38316; b = 18392; cin = 0;
#10 a = 54287; b = 39786; cin = 0;
#10 a = 10918; b = 17723; cin = 0;
#10 a = 69135; b = 25870; cin = 0;
#10 a = 56543; b = 49431; cin = 0;
#10 a = 24499; b = 41435; cin = 1;
#10 a = 25096; b = 62306; cin = 0;
#10 a = 40069; b = 15447; cin = 1;
#10 a = 53138; b = 22630; cin = 1;
#10 a = 62851; b = 59225; cin = 0;
#10 a = 69978; b = 27541; cin = 0;
#10 a = 51947; b = 58180; cin = 0;
#10 a = 17785; b = 69098; cin = 1;
#10 a = 24992; b = 68233; cin = 0;
#10 a = 782; b = 31128; cin = 1;
#10 a = 15130; b = 55627; cin = 0;
#10 a = 31170; b = 57076; cin = 1;
#10 a = 54472; b = 27145; cin = 0;
#10 a = 20925; b = 10283; cin = 1;
#10 a = 11397; b = 49486; cin = 0;
#10 a = 51863; b = 25817; cin = 1;
#10 a = 40721; b = 54116; cin = 0;
#10 a = 69365; b = 48253; cin = 0;
#10 a = 22085; b = 3245; cin = 0;
#10 a = 675; b = 4027; cin = 0;
#10 a = 5048; b = 65510; cin = 0;
#10 a = 3560; b = 26680; cin = 0;
#10 a = 18027; b = 57504; cin = 1;
#10 a = 646; b = 8430; cin = 0;
#10 a = 29543; b = 66179; cin = 1;
#10 a = 24017; b = 48042; cin = 0;
#10 a = 46032; b = 65115; cin = 0;
#10 a = 32580; b = 40832; cin = 1;
#10 a = 64579; b = 62917; cin = 1;
#10 a = 1163; b = 63592; cin = 0;
#10 a = 38875; b = 44992; cin = 0;
#10 a = 62215; b = 24905; cin = 0;
#10 a = 2631; b = 42932; cin = 1;
#10 a = 16544; b = 43578; cin = 1;
#10 a = 17093; b = 49473; cin = 0;
#10 a = 67128; b = 3490; cin = 0;
#10 a = 2980; b = 49523; cin = 1;
#10 a = 62948; b = 58455; cin = 1;
#10 a = 7521; b = 29386; cin = 1;
#10 a = 48988; b = 30549; cin = 1;
#10 a = 47187; b = 69425; cin = 0;
#10 a = 40895; b = 37992; cin = 1;
#10 a = 37636; b = 40624; cin = 1;
#10 a = 68233; b = 33520; cin = 0;
#10 a = 37260; b = 50613; cin = 1;
#10 a = 2466; b = 47741; cin = 0;
#10 a = 62066; b = 50721; cin = 1;
#10 a = 46781; b = 20021; cin = 0;
#10 a = 48680; b = 27543; cin = 1;
#10 a = 67145; b = 52883; cin = 0;
#10 a = 31907; b = 30070; cin = 1;
#10 a = 18013; b = 966; cin = 0;
#10 a = 52672; b = 14954; cin = 0;
#10 a = 12967; b = 13187; cin = 0;
#10 a = 16841; b = 50447; cin = 0;
#10 a = 189; b = 52913; cin = 1;
#10 a = 33379; b = 21331; cin = 1;
#10 a = 46092; b = 44464; cin = 0;
#10 a = 23612; b = 23144; cin = 1;
#10 a = 6871; b = 66642; cin = 1;
#10 a = 44328; b = 28549; cin = 1;
#10 a = 33913; b = 46562; cin = 1;
#10 a = 15139; b = 5586; cin = 1;
#10 a = 59693; b = 64905; cin = 0;
#10 a = 67768; b = 11747; cin = 1;
#10 a = 56456; b = 58288; cin = 0;
#10 a = 69237; b = 21667; cin = 1;
#10 a = 39092; b = 44111; cin = 1;
#10 a = 28969; b = 44075; cin = 0;
#10 a = 22740; b = 50947; cin = 0;
#10 a = 69395; b = 1627; cin = 1;
#10 a = 6121; b = 35540; cin = 1;
#10 a = 36516; b = 27032; cin = 1;
#10 a = 35514; b = 16725; cin = 0;
#10 a = 24050; b = 14493; cin = 1;
#10 a = 39386; b = 47301; cin = 1;
#10 a = 37634; b = 46539; cin = 0;
#10 a = 33566; b = 15631; cin = 1;
#10 a = 50313; b = 20952; cin = 1;
#10 a = 43853; b = 43693; cin = 0;
#10 a = 10387; b = 43088; cin = 1;
#10 a = 51822; b = 25561; cin = 1;
#10 a = 46171; b = 62078; cin = 1;
#10 a = 22458; b = 3944; cin = 1;
#10 a = 17299; b = 27994; cin = 0;
#10 a = 238; b = 43732; cin = 0;
#10 a = 17818; b = 57719; cin = 1;
#10 a = 57064; b = 67637; cin = 0;
#10 a = 46774; b = 47950; cin = 1;
#10 a = 10559; b = 68156; cin = 0;
#10 a = 1643; b = 54895; cin = 0;
#10 a = 64354; b = 36718; cin = 0;
#10 a = 68957; b = 59241; cin = 0;
#10 a = 30593; b = 11700; cin = 0;
#10 a = 8954; b = 5351; cin = 0;
#10 a = 48160; b = 51941; cin = 1;
#10 a = 41020; b = 69759; cin = 0;
#10 a = 10419; b = 56824; cin = 1;
#10 a = 18154; b = 9950; cin = 1;
#10 a = 489; b = 20509; cin = 1;
#10 a = 26517; b = 22152; cin = 1;
#10 a = 1985; b = 62858; cin = 1;
#10 a = 3015; b = 61815; cin = 0;
#10 a = 42475; b = 22408; cin = 0;
#10 a = 39527; b = 31362; cin = 1;
#10 a = 17278; b = 55875; cin = 1;
#10 a = 38761; b = 3247; cin = 0;
#10 a = 47963; b = 13667; cin = 0;
#10 a = 31154; b = 31821; cin = 0;
#10 a = 62295; b = 8662; cin = 1;
#10 a = 21593; b = 11531; cin = 1;
#10 a = 12138; b = 59868; cin = 1;
#10 a = 39401; b = 39236; cin = 1;
#10 a = 55905; b = 11711; cin = 1;
#10 a = 14110; b = 27591; cin = 0;
#10 a = 24017; b = 44869; cin = 1;
#10 a = 15866; b = 13630; cin = 0;
#10 a = 7475; b = 37945; cin = 1;
#10 a = 8611; b = 69099; cin = 0;
#10 a = 43346; b = 61394; cin = 0;
#10 a = 4941; b = 59339; cin = 1;
#10 a = 58689; b = 1477; cin = 0;
#10 a = 11646; b = 40878; cin = 0;
#10 a = 50067; b = 26784; cin = 1;
#10 a = 17249; b = 17246; cin = 0;
#10 a = 62145; b = 17615; cin = 1;
#10 a = 22916; b = 33482; cin = 1;
#10 a = 33286; b = 17309; cin = 0;
#10 a = 57324; b = 25920; cin = 1;
#10 a = 19534; b = 45618; cin = 0;
#10 a = 60407; b = 26912; cin = 1;
#10 a = 19162; b = 15601; cin = 1;
#10 a = 37786; b = 3599; cin = 1;
#10 a = 25646; b = 53667; cin = 1;
#10 a = 25218; b = 47268; cin = 1;
#10 a = 52380; b = 39413; cin = 1;
#10 a = 30764; b = 38681; cin = 1;
#10 a = 22777; b = 1967; cin = 0;
#10 a = 29088; b = 35643; cin = 0;
#10 a = 34497; b = 55178; cin = 1;
#10 a = 54005; b = 21937; cin = 1;
#10 a = 16501; b = 41099; cin = 0;
#10 a = 3178; b = 55238; cin = 1;
#10 a = 30733; b = 10884; cin = 0;
#10 a = 61425; b = 36102; cin = 0;
#10 a = 15714; b = 64835; cin = 1;
#10 a = 57619; b = 25599; cin = 0;
#10 a = 39358; b = 24728; cin = 0;
#10 a = 14758; b = 30168; cin = 1;
#10 a = 62431; b = 41018; cin = 1;
#10 a = 15722; b = 25023; cin = 0;
#10 a = 65925; b = 17876; cin = 0;
#10 a = 38081; b = 21054; cin = 0;
#10 a = 37484; b = 28140; cin = 0;
#10 a = 43259; b = 65917; cin = 1;
#10 a = 26301; b = 11631; cin = 0;
#10 a = 25109; b = 45603; cin = 1;
#10 a = 38949; b = 61313; cin = 1;
#10 a = 31109; b = 52424; cin = 0;
#10 a = 12561; b = 44855; cin = 0;
#10 a = 25542; b = 60577; cin = 1;
#10 a = 36813; b = 56502; cin = 0;
#10 a = 19183; b = 24583; cin = 0;
#10 a = 33143; b = 38419; cin = 0;
#10 a = 34339; b = 58030; cin = 1;
#10 a = 1638; b = 14332; cin = 1;
#10 a = 10124; b = 15793; cin = 0;
#10 a = 20561; b = 31094; cin = 1;
#10 a = 32079; b = 62204; cin = 1;
#10 a = 3765; b = 51117; cin = 0;
#10 a = 16469; b = 53011; cin = 1;
#10 a = 54196; b = 19824; cin = 1;
#10 a = 16152; b = 15359; cin = 0;
#10 a = 69163; b = 24854; cin = 0;
#10 a = 10313; b = 59194; cin = 0;
#10 a = 17381; b = 60832; cin = 0;
#10 a = 12432; b = 47309; cin = 1;
#10 a = 29438; b = 67870; cin = 0;
#10 a = 14109; b = 29949; cin = 0;
#10 a = 4853; b = 10066; cin = 1;
#10 a = 16803; b = 26535; cin = 0;
#10 a = 65683; b = 57084; cin = 1;
#10 a = 31064; b = 3236; cin = 0;
#10 a = 67381; b = 2399; cin = 1;
#10 a = 2117; b = 59065; cin = 1;
#10 a = 64883; b = 6446; cin = 1;
#10 a = 48334; b = 65230; cin = 0;
#10 a = 23929; b = 1020; cin = 1;
#10 a = 6971; b = 15129; cin = 0;
#10 a = 52217; b = 66334; cin = 1;
#10 a = 54932; b = 59490; cin = 0;
#10 a = 40659; b = 55173; cin = 0;
#10 a = 22562; b = 62589; cin = 1;
#10 a = 66176; b = 59970; cin = 0;
#10 a = 64645; b = 62087; cin = 1;
#10 a = 28660; b = 33323; cin = 1;
#10 a = 53508; b = 58009; cin = 1;
#10 a = 32016; b = 58290; cin = 1;
#10 a = 54747; b = 65262; cin = 1;
#10 a = 37428; b = 23831; cin = 1;
#10 a = 30175; b = 8764; cin = 1;
#10 a = 25809; b = 25775; cin = 0;
#10 a = 54880; b = 24689; cin = 0;
#10 a = 40835; b = 20865; cin = 0;
#10 a = 51893; b = 61863; cin = 0;
#10 a = 52017; b = 66875; cin = 1;
#10 a = 58586; b = 50383; cin = 0;
#10 a = 13090; b = 58752; cin = 0;
#10 a = 62261; b = 43499; cin = 0;
#10 a = 32914; b = 10927; cin = 0;
#10 a = 69902; b = 17454; cin = 0;
#10 a = 26379; b = 19616; cin = 1;
#10 a = 14382; b = 50848; cin = 0;
#10 a = 64974; b = 21683; cin = 1;
#10 a = 35536; b = 49928; cin = 0;
#10 a = 44538; b = 31945; cin = 0;
#10 a = 63215; b = 66884; cin = 1;
#10 a = 69901; b = 9974; cin = 1;
#10 a = 64878; b = 48587; cin = 1;
#10 a = 55116; b = 57854; cin = 0;
#10 a = 45538; b = 57756; cin = 1;
#10 a = 44724; b = 60487; cin = 1;
#10 a = 69685; b = 4869; cin = 1;
#10 a = 25687; b = 69843; cin = 0;
#10 a = 48907; b = 35380; cin = 0;
#10 a = 40341; b = 56270; cin = 0;
#10 a = 52299; b = 49486; cin = 0;
#10 a = 20993; b = 25739; cin = 0;
#10 a = 24790; b = 20617; cin = 1;
#10 a = 2087; b = 52086; cin = 1;
#10 a = 36664; b = 27624; cin = 1;
#10 a = 65047; b = 2349; cin = 1;
#10 a = 43046; b = 48386; cin = 0;
#10 a = 48245; b = 50426; cin = 0;
#10 a = 5127; b = 29333; cin = 0;
#10 a = 58289; b = 69674; cin = 0;
#10 a = 49749; b = 28326; cin = 0;
#10 a = 38093; b = 25671; cin = 0;
#10 a = 12763; b = 50461; cin = 1;
#10 a = 12373; b = 28901; cin = 1;
#10 a = 69836; b = 65565; cin = 0;
#10 a = 45056; b = 36964; cin = 1;
#10 a = 57115; b = 10010; cin = 1;
#10 a = 50395; b = 34607; cin = 1;
#10 a = 43519; b = 16086; cin = 0;
#10 a = 2023; b = 50727; cin = 1;
#10 a = 39502; b = 30477; cin = 1;
#10 a = 56466; b = 44922; cin = 0;
#10 a = 29170; b = 57686; cin = 1;
#10 a = 68844; b = 59; cin = 0;
#10 a = 20603; b = 69895; cin = 1;
#10 a = 69987; b = 21303; cin = 1;
#10 a = 28072; b = 54770; cin = 1;
#10 a = 10896; b = 35166; cin = 0;
#10 a = 67793; b = 8685; cin = 0;
#10 a = 60376; b = 57061; cin = 0;
#10 a = 28985; b = 26563; cin = 1;
#10 a = 2272; b = 59381; cin = 1;
#10 a = 24878; b = 64904; cin = 1;
#10 a = 50649; b = 40100; cin = 0;
#10 a = 11674; b = 60703; cin = 0;
#10 a = 38263; b = 37043; cin = 1;
#10 a = 31817; b = 41467; cin = 0;
#10 a = 58084; b = 52363; cin = 0;
#10 a = 48959; b = 26509; cin = 1;
#10 a = 55919; b = 63237; cin = 0;
#10 a = 43607; b = 22222; cin = 1;
#10 a = 38124; b = 846; cin = 1;
#10 a = 7564; b = 25724; cin = 1;
#10 a = 11041; b = 52725; cin = 1;
#10 a = 14578; b = 64399; cin = 0;
#10 a = 64362; b = 9015; cin = 1;
#10 a = 41801; b = 40832; cin = 1;
#10 a = 4011; b = 5268; cin = 0;
#10 a = 24091; b = 54227; cin = 1;
#10 a = 52857; b = 40147; cin = 0;
#10 a = 45035; b = 60106; cin = 0;
#10 a = 40129; b = 28231; cin = 0;
#10 a = 956; b = 12147; cin = 0;
#10 a = 50335; b = 23188; cin = 0;
#10 a = 46166; b = 14118; cin = 1;
#10 a = 9052; b = 8480; cin = 0;
#10 a = 8982; b = 26634; cin = 0;
#10 a = 26731; b = 6997; cin = 1;
#10 a = 3195; b = 31089; cin = 0;
#10 a = 6169; b = 60298; cin = 1;
#10 a = 2379; b = 11685; cin = 0;
#10 a = 67164; b = 51814; cin = 1;
#10 a = 62794; b = 29122; cin = 0;
#10 a = 60501; b = 9457; cin = 0;
#10 a = 40933; b = 31975; cin = 1;
#10 a = 38468; b = 41028; cin = 1;
#10 a = 68667; b = 26362; cin = 1;
#10 a = 46049; b = 53093; cin = 1;
#10 a = 5052; b = 56288; cin = 0;
#10 a = 41931; b = 62457; cin = 0;
#10 a = 25308; b = 41189; cin = 1;
#10 a = 45144; b = 38353; cin = 0;
#10 a = 23211; b = 31147; cin = 0;
#10 a = 59777; b = 21648; cin = 0;
#10 a = 25884; b = 38933; cin = 1;
#10 a = 6109; b = 7402; cin = 1;
#10 a = 41166; b = 52421; cin = 1;
#10 a = 9210; b = 4822; cin = 0;
#10 a = 54251; b = 9875; cin = 1;
#10 a = 36733; b = 28158; cin = 0;
#10 a = 9513; b = 29818; cin = 1;
#10 a = 63978; b = 4963; cin = 0;
#10 a = 6610; b = 28174; cin = 0;
#10 a = 48365; b = 64304; cin = 0;
#10 a = 52281; b = 20188; cin = 0;
#10 a = 41820; b = 2649; cin = 0;
#10 a = 25092; b = 20167; cin = 1;
#10 a = 58373; b = 29377; cin = 1;
#10 a = 27452; b = 59980; cin = 0;
#10 a = 52819; b = 26713; cin = 0;
#10 a = 643; b = 12578; cin = 1;
#10 a = 36009; b = 6557; cin = 0;
#10 a = 39727; b = 59519; cin = 0;
#10 a = 50945; b = 14236; cin = 0;
#10 a = 13812; b = 66517; cin = 0;
#10 a = 61964; b = 14690; cin = 1;
#10 a = 47518; b = 39782; cin = 1;
#10 a = 61845; b = 4507; cin = 0;
#10 a = 10994; b = 31959; cin = 1;
#10 a = 40019; b = 14778; cin = 0;
#10 a = 27201; b = 61774; cin = 1;
#10 a = 20554; b = 4135; cin = 0;
#10 a = 18870; b = 43862; cin = 1;
#10 a = 21713; b = 1160; cin = 0;
#10 a = 18859; b = 14972; cin = 1;
#10 a = 12546; b = 6936; cin = 1;
#10 a = 8881; b = 30806; cin = 1;
#10 a = 1736; b = 22651; cin = 1;
#10 a = 23969; b = 33645; cin = 0;
#10 a = 36182; b = 50016; cin = 1;
#10 a = 51460; b = 53570; cin = 1;
#10 a = 9317; b = 4124; cin = 0;
#10 a = 20083; b = 69347; cin = 0;
#10 a = 66721; b = 67412; cin = 0;
#10 a = 57595; b = 16271; cin = 0;
#10 a = 21338; b = 5169; cin = 0;
#10 a = 69772; b = 60403; cin = 0;
#10 a = 17987; b = 62139; cin = 1;
#10 a = 17062; b = 16108; cin = 1;
#10 a = 48097; b = 28642; cin = 1;
#10 a = 23910; b = 56455; cin = 1;
#10 a = 37849; b = 42124; cin = 0;
#10 a = 55923; b = 38560; cin = 1;
#10 a = 47859; b = 35281; cin = 1;
#10 a = 17308; b = 69228; cin = 0;
#10 a = 48080; b = 20566; cin = 0;
#10 a = 15789; b = 20338; cin = 1;
#10 a = 60655; b = 14678; cin = 0;
#10 a = 34525; b = 31740; cin = 1;
#10 a = 18392; b = 9837; cin = 1;
#10 a = 28627; b = 10099; cin = 0;
#10 a = 46081; b = 47948; cin = 1;
#10 a = 20363; b = 33871; cin = 1;
#10 a = 63992; b = 58083; cin = 0;
#10 a = 35033; b = 5391; cin = 0;
#10 a = 68697; b = 29823; cin = 0;
#10 a = 37531; b = 45612; cin = 1;
#10 a = 43120; b = 12620; cin = 1;
#10 a = 64497; b = 23497; cin = 1;
#10 a = 54686; b = 18241; cin = 1;
#10 a = 3517; b = 46868; cin = 0;
#10 a = 8804; b = 69301; cin = 1;
#10 a = 56215; b = 66016; cin = 0;
#10 a = 2186; b = 60008; cin = 1;
#10 a = 29790; b = 1393; cin = 0;
#10 a = 56622; b = 46443; cin = 0;
#10 a = 10372; b = 13974; cin = 0;
#10 a = 30813; b = 33447; cin = 0;
#10 a = 42284; b = 27944; cin = 1;
#10 a = 15496; b = 58982; cin = 0;
#10 a = 44897; b = 62499; cin = 1;
#10 a = 60749; b = 1303; cin = 0;
#10 a = 8198; b = 57518; cin = 1;
#10 a = 35871; b = 59704; cin = 1;
#10 a = 27978; b = 65846; cin = 1;
#10 a = 25477; b = 52468; cin = 0;
#10 a = 52799; b = 39193; cin = 0;
#10 a = 32085; b = 46358; cin = 1;
#10 a = 344; b = 18643; cin = 1;
#10 a = 38451; b = 10491; cin = 1;
#10 a = 1152; b = 31740; cin = 1;
#10 a = 10721; b = 22489; cin = 0;
#10 a = 65943; b = 7040; cin = 1;
#10 a = 23534; b = 42911; cin = 1;
#10 a = 41134; b = 47241; cin = 0;
#10 a = 36479; b = 2718; cin = 0;
#10 a = 8267; b = 31869; cin = 1;
#10 a = 40381; b = 40307; cin = 0;
#10 a = 35943; b = 40651; cin = 1;
#10 a = 35800; b = 55454; cin = 0;
#10 a = 992; b = 56606; cin = 0;
#10 a = 52331; b = 43679; cin = 1;
#10 a = 11325; b = 15975; cin = 1;
#10 a = 27838; b = 39509; cin = 0;
#10 a = 10408; b = 10643; cin = 0;
#10 a = 58824; b = 23474; cin = 0;
#10 a = 19708; b = 8093; cin = 0;
#10 a = 66138; b = 48475; cin = 1;
#10 a = 18926; b = 60770; cin = 0;
#10 a = 36709; b = 2922; cin = 0;
#10 a = 64983; b = 3914; cin = 1;
#10 a = 54997; b = 32597; cin = 0;
#10 a = 67500; b = 43923; cin = 1;
#10 a = 17044; b = 1761; cin = 1;
#10 a = 55850; b = 12169; cin = 0;
#10 a = 1898; b = 993; cin = 1;
#10 a = 67017; b = 67054; cin = 0;
#10 a = 357; b = 63192; cin = 1;
#10 a = 67652; b = 58470; cin = 1;
#10 a = 11950; b = 25179; cin = 0;
#10 a = 58054; b = 20162; cin = 0;
#10 a = 67117; b = 5159; cin = 0;
#10 a = 49860; b = 2659; cin = 1;
#10 a = 48577; b = 66055; cin = 0;
#10 a = 16804; b = 51906; cin = 0;
#10 a = 18379; b = 30156; cin = 1;
#10 a = 43428; b = 3525; cin = 1;
#10 a = 6570; b = 3882; cin = 1;
#10 a = 18188; b = 1534; cin = 1;
#10 a = 43279; b = 59836; cin = 0;
#10 a = 1293; b = 24243; cin = 0;
#10 a = 9574; b = 21360; cin = 1;
#10 a = 50452; b = 47572; cin = 1;
#10 a = 18901; b = 26150; cin = 0;
#10 a = 11815; b = 19306; cin = 0;
#10 a = 40547; b = 37685; cin = 1;
#10 a = 22977; b = 57465; cin = 0;
#10 a = 26108; b = 64036; cin = 1;
#10 a = 68784; b = 58576; cin = 1;
#10 a = 29929; b = 31855; cin = 0;
#10 a = 62606; b = 9501; cin = 1;
#10 a = 21796; b = 19075; cin = 1;
#10 a = 56146; b = 69527; cin = 0;
#10 a = 23155; b = 64780; cin = 0;
#10 a = 8923; b = 6595; cin = 0;
#10 a = 246; b = 23495; cin = 0;
#10 a = 44429; b = 46472; cin = 1;
#10 a = 22137; b = 48932; cin = 1;
#10 a = 50080; b = 24068; cin = 1;
#10 a = 9558; b = 53998; cin = 1;
#10 a = 51576; b = 22956; cin = 0;
#10 a = 1485; b = 44752; cin = 1;
#10 a = 19106; b = 30898; cin = 0;
#10 a = 60652; b = 30405; cin = 0;
#10 a = 58348; b = 39329; cin = 1;
#10 a = 5351; b = 15927; cin = 0;
#10 a = 12743; b = 36708; cin = 0;
#10 a = 31248; b = 58845; cin = 1;
#10 a = 20142; b = 38926; cin = 1;
#10 a = 67611; b = 24836; cin = 1;
#10 a = 6936; b = 6412; cin = 1;
#10 a = 2114; b = 54249; cin = 0;
#10 a = 16367; b = 49707; cin = 0;
#10 a = 30147; b = 40360; cin = 0;
#10 a = 15059; b = 28708; cin = 1;
#10 a = 52919; b = 10411; cin = 0;
#10 a = 44273; b = 23154; cin = 0;
#10 a = 58452; b = 30755; cin = 1;
#10 a = 51563; b = 50897; cin = 1;
#10 a = 68742; b = 48508; cin = 1;
#10 a = 46272; b = 31797; cin = 1;
#10 a = 23109; b = 33911; cin = 0;
#10 a = 21051; b = 50279; cin = 0;
#10 a = 49892; b = 56778; cin = 0;
#10 a = 39138; b = 48190; cin = 0;
#10 a = 20417; b = 31109; cin = 0;
#10 a = 17623; b = 5382; cin = 0;
#10 a = 51537; b = 63834; cin = 1;
#10 a = 50648; b = 21749; cin = 0;
#10 a = 18686; b = 20492; cin = 1;
#10 a = 34263; b = 43116; cin = 0;
#10 a = 56253; b = 42577; cin = 1;
#10 a = 38843; b = 63629; cin = 0;
#10 a = 47493; b = 43521; cin = 1;
#10 a = 26503; b = 59011; cin = 1;
#10 a = 10574; b = 55780; cin = 0;
#10 a = 5056; b = 3403; cin = 0;
#10 a = 69044; b = 54940; cin = 1;
#10 a = 23788; b = 35588; cin = 0;
#10 a = 29428; b = 30626; cin = 0;
#10 a = 59929; b = 64890; cin = 0;
#10 a = 28579; b = 27495; cin = 0;
#10 a = 7493; b = 42690; cin = 1;
#10 a = 13037; b = 20184; cin = 0;
#10 a = 5360; b = 46687; cin = 1;
#10 a = 22225; b = 33613; cin = 1;
#10 a = 199; b = 38669; cin = 0;
#10 a = 53556; b = 14066; cin = 0;
#10 a = 53451; b = 37854; cin = 0;
#10 a = 28743; b = 67282; cin = 1;
#10 a = 880; b = 33564; cin = 1;
#10 a = 62484; b = 38495; cin = 0;
#10 a = 3018; b = 45988; cin = 0;
#10 a = 7181; b = 59026; cin = 0;
#10 a = 31217; b = 40738; cin = 0;
#10 a = 44264; b = 62964; cin = 1;
#10 a = 19443; b = 39515; cin = 1;
#10 a = 68025; b = 69423; cin = 1;
#10 a = 7899; b = 52874; cin = 1;
#10 a = 29714; b = 57970; cin = 1;
#10 a = 58507; b = 35202; cin = 1;
#10 a = 12190; b = 27686; cin = 1;
#10 a = 39720; b = 7057; cin = 1;
#10 a = 63588; b = 14238; cin = 1;
#10 a = 60345; b = 45456; cin = 0;
#10 a = 33789; b = 66072; cin = 0;
#10 a = 40846; b = 15516; cin = 1;
#10 a = 62925; b = 59893; cin = 1;
#10 a = 5422; b = 67793; cin = 1;
#10 a = 55773; b = 3859; cin = 1;
#10 a = 33407; b = 62366; cin = 1;
#10 a = 20956; b = 50908; cin = 0;
#10 a = 47001; b = 20628; cin = 1;
#10 a = 25387; b = 60568; cin = 1;
#10 a = 39150; b = 50913; cin = 1;
#10 a = 23652; b = 14702; cin = 0;
#10 a = 47470; b = 55549; cin = 0;
#10 a = 17156; b = 24826; cin = 1;
#10 a = 9913; b = 6601; cin = 0;
#10 a = 31896; b = 62374; cin = 1;
#10 a = 41850; b = 2133; cin = 1;
#10 a = 17005; b = 69442; cin = 1;
#10 a = 66199; b = 22795; cin = 1;
#10 a = 52450; b = 48182; cin = 0;
#10 a = 52940; b = 63685; cin = 1;
#10 a = 5237; b = 17337; cin = 0;
#10 a = 23607; b = 41160; cin = 1;
#10 a = 33845; b = 34668; cin = 1;
#10 a = 33977; b = 44581; cin = 0;
#10 a = 31901; b = 52829; cin = 1;
#10 a = 56389; b = 1031; cin = 0;
#10 a = 3242; b = 18037; cin = 0;
#10 a = 1004; b = 60588; cin = 0;
#10 a = 19393; b = 43039; cin = 0;
#10 a = 4703; b = 2331; cin = 1;
#10 a = 64575; b = 53920; cin = 1;
#10 a = 21853; b = 53880; cin = 1;
#10 a = 34680; b = 17725; cin = 1;
#10 a = 48685; b = 51702; cin = 0;
#10 a = 45644; b = 59956; cin = 1;
#10 a = 34977; b = 46345; cin = 1;
#10 a = 2795; b = 49587; cin = 0;
#10 a = 40056; b = 50591; cin = 0;
#10 a = 30112; b = 46337; cin = 1;
#10 a = 44702; b = 51040; cin = 0;
#10 a = 52978; b = 21967; cin = 1;
#10 a = 31295; b = 43820; cin = 1;
#10 a = 50772; b = 54852; cin = 0;
#10 a = 34917; b = 33538; cin = 1;
#10 a = 39995; b = 55534; cin = 1;
#10 a = 27902; b = 20511; cin = 0;
#10 a = 63193; b = 23306; cin = 1;
#10 a = 46521; b = 39714; cin = 1;
#10 a = 66790; b = 69826; cin = 0;
#10 a = 36449; b = 20881; cin = 0;
#10 a = 54792; b = 50211; cin = 0;
#10 a = 57055; b = 11506; cin = 0;
#10 a = 43198; b = 62278; cin = 1;
#10 a = 23418; b = 27195; cin = 1;
#10 a = 55341; b = 43542; cin = 1;
#10 a = 53572; b = 1444; cin = 0;
#10 a = 4500; b = 40990; cin = 0;
#10 a = 5016; b = 63863; cin = 1;
#10 a = 32475; b = 37005; cin = 1;
#10 a = 36271; b = 3455; cin = 0;
#10 a = 67459; b = 58247; cin = 1;
#10 a = 26967; b = 45302; cin = 1;
#10 a = 30296; b = 64852; cin = 1;
#10 a = 18477; b = 18270; cin = 0;
#10 a = 16548; b = 3612; cin = 0;
#10 a = 46505; b = 33536; cin = 1;
#10 a = 50621; b = 38037; cin = 1;
#10 a = 30747; b = 19405; cin = 0;
#10 a = 50588; b = 51880; cin = 0;
#10 a = 46608; b = 64503; cin = 1;
#10 a = 63508; b = 61962; cin = 0;
#10 a = 36972; b = 18930; cin = 0;
#10 a = 21941; b = 25578; cin = 0;
#10 a = 45541; b = 44055; cin = 0;
#10 a = 2687; b = 36955; cin = 0;
#10 a = 27024; b = 13460; cin = 1;
#10 a = 5509; b = 40433; cin = 0;
#10 a = 24984; b = 47532; cin = 1;
#10 a = 38322; b = 28121; cin = 1;
#10 a = 18666; b = 4729; cin = 0;
#10 a = 2465; b = 68237; cin = 0;
#10 a = 67215; b = 11561; cin = 0;
#10 a = 37267; b = 33503; cin = 0;
#10 a = 2171; b = 55396; cin = 1;
#10 a = 31698; b = 58083; cin = 0;
#10 a = 64836; b = 61459; cin = 0;
#10 a = 37863; b = 66968; cin = 1;
#10 a = 25279; b = 21952; cin = 0;
#10 a = 55748; b = 36627; cin = 1;
#10 a = 44449; b = 55293; cin = 0;
#10 a = 4005; b = 34111; cin = 1;
#10 a = 25524; b = 31326; cin = 1;
#10 a = 65972; b = 68594; cin = 0;
#10 a = 38351; b = 47117; cin = 0;
#10 a = 31136; b = 8815; cin = 1;
#10 a = 37229; b = 50004; cin = 1;
#10 a = 56781; b = 17867; cin = 1;
#10 a = 23119; b = 43147; cin = 0;
#10 a = 36989; b = 5247; cin = 1;
#10 a = 55332; b = 26049; cin = 0;
#10 a = 8404; b = 30054; cin = 1;
#10 a = 29713; b = 55578; cin = 0;
#10 a = 38936; b = 27903; cin = 0;
#10 a = 58014; b = 42606; cin = 1;
#10 a = 62488; b = 50094; cin = 1;
#10 a = 55046; b = 17323; cin = 1;
#10 a = 15415; b = 4105; cin = 0;
#10 a = 19104; b = 3576; cin = 1;
#10 a = 44746; b = 40565; cin = 1;
#10 a = 13367; b = 25897; cin = 0;
#10 a = 60930; b = 34301; cin = 0;
#10 a = 48955; b = 40366; cin = 1;
#10 a = 44659; b = 55655; cin = 0;
#10 a = 38957; b = 20021; cin = 0;
#10 a = 56725; b = 12510; cin = 0;
#10 a = 59660; b = 43908; cin = 0;
#10 a = 42599; b = 35675; cin = 1;
#10 a = 43405; b = 54779; cin = 1;
#10 a = 17359; b = 5878; cin = 0;
#10 a = 19264; b = 19245; cin = 1;
#10 a = 866; b = 56527; cin = 0;
#10 a = 12522; b = 11835; cin = 0;
#10 a = 56109; b = 56494; cin = 1;
#10 a = 33951; b = 1804; cin = 1;
#10 a = 8047; b = 34881; cin = 1;
#10 a = 8590; b = 24541; cin = 1;
#10 a = 26456; b = 67140; cin = 0;
#10 a = 24779; b = 16897; cin = 1;
#10 a = 26678; b = 34256; cin = 1;
#10 a = 45494; b = 53520; cin = 1;
#10 a = 66559; b = 30738; cin = 0;
#10 a = 28277; b = 19613; cin = 1;
#10 a = 6713; b = 5722; cin = 0;
#10 a = 40805; b = 16026; cin = 0;
#10 a = 1270; b = 24073; cin = 1;
#10 a = 44245; b = 9015; cin = 0;
#10 a = 37480; b = 35471; cin = 0;
#10 a = 20038; b = 36602; cin = 1;
#10 a = 33727; b = 63280; cin = 0;
#10 a = 53295; b = 15126; cin = 0;
#10 a = 22108; b = 11685; cin = 1;
#10 a = 47448; b = 39962; cin = 0;
#10 a = 60976; b = 46676; cin = 0;
#10 a = 60998; b = 63833; cin = 0;
#10 a = 39176; b = 65103; cin = 0;
#10 a = 5883; b = 15700; cin = 1;
#10 a = 19835; b = 53180; cin = 1;
#10 a = 30927; b = 3218; cin = 1;
#10 a = 35268; b = 13297; cin = 0;
#10 a = 3866; b = 42944; cin = 0;
#10 a = 2337; b = 65052; cin = 0;
#10 a = 31546; b = 18853; cin = 0;
#10 a = 56720; b = 56181; cin = 0;
#10 a = 63968; b = 47179; cin = 1;
#10 a = 17243; b = 16355; cin = 0;
#10 a = 64591; b = 68590; cin = 0;
#10 a = 27306; b = 64777; cin = 0;
#10 a = 25493; b = 25704; cin = 0;
#10 a = 36635; b = 60972; cin = 0;
#10 a = 41057; b = 41191; cin = 0;
#10 a = 60605; b = 43528; cin = 1;
#10 a = 21839; b = 51426; cin = 0;
#10 a = 69388; b = 14498; cin = 1;
#10 a = 46316; b = 8466; cin = 0;
#10 a = 40726; b = 25709; cin = 1;
#10 a = 52942; b = 66652; cin = 1;
#10 a = 10859; b = 23959; cin = 0;
#10 a = 21955; b = 25804; cin = 0;
#10 a = 12622; b = 62439; cin = 0;
#10 a = 16586; b = 33496; cin = 1;
#10 a = 39846; b = 24102; cin = 1;
#10 a = 58159; b = 45941; cin = 1;
#10 a = 1677; b = 21681; cin = 1;
#10 a = 1376; b = 67998; cin = 0;
#10 a = 24606; b = 15076; cin = 1;
#10 a = 40543; b = 44370; cin = 0;
#10 a = 31422; b = 55229; cin = 1;
#10 a = 40726; b = 7185; cin = 1;
#10 a = 52086; b = 19807; cin = 1;
#10 a = 30771; b = 12745; cin = 1;
#10 a = 26998; b = 52591; cin = 1;
#10 a = 20402; b = 17103; cin = 1;
#10 a = 17935; b = 65132; cin = 0;
#10 a = 53615; b = 42861; cin = 0;
#10 a = 4113; b = 43819; cin = 0;
#10 a = 26672; b = 14363; cin = 1;
#10 a = 69532; b = 45785; cin = 0;
#10 a = 19055; b = 62864; cin = 1;
#10 a = 18031; b = 21302; cin = 0;
#10 a = 9446; b = 28425; cin = 1;
#10 a = 34357; b = 55424; cin = 1;
#10 a = 13371; b = 52178; cin = 0;
#10 a = 61030; b = 113; cin = 0;
#10 a = 60370; b = 53728; cin = 1;
#10 a = 34061; b = 34193; cin = 1;
#10 a = 69179; b = 60866; cin = 0;
#10 a = 8668; b = 36750; cin = 1;
#10 a = 3387; b = 55806; cin = 1;
#10 a = 27994; b = 3837; cin = 0;
#10 a = 2409; b = 59635; cin = 1;
#10 a = 35920; b = 23992; cin = 1;
#10 a = 52023; b = 13715; cin = 1;
#10 a = 61581; b = 4745; cin = 1;
#10 a = 66272; b = 41468; cin = 1;
#10 a = 43823; b = 5529; cin = 1;
#10 a = 41546; b = 4708; cin = 1;
#10 a = 53632; b = 13377; cin = 1;
#10 a = 17856; b = 63116; cin = 1;
#10 a = 21295; b = 21110; cin = 0;
#10 a = 69685; b = 69871; cin = 1;
#10 a = 6501; b = 35792; cin = 0;
#10 a = 45092; b = 64167; cin = 1;
#10 a = 65862; b = 55749; cin = 1;
#10 a = 16745; b = 52021; cin = 1;
#10 a = 21356; b = 2196; cin = 0;
#10 a = 12865; b = 20095; cin = 0;
#10 a = 65240; b = 3727; cin = 1;
#10 a = 60718; b = 67935; cin = 1;
#10 a = 18353; b = 19231; cin = 0;
#10 a = 26178; b = 65268; cin = 1;
#10 a = 23637; b = 1769; cin = 1;
#10 a = 45089; b = 23214; cin = 1;
#10 a = 32961; b = 19076; cin = 0;
#10 a = 25578; b = 35821; cin = 1;
#10 a = 36015; b = 33529; cin = 1;
#10 a = 5629; b = 46395; cin = 0;
#10 a = 26303; b = 17987; cin = 0;
#10 a = 36707; b = 8705; cin = 1;
#10 a = 40226; b = 3411; cin = 0;
#10 a = 41208; b = 29589; cin = 1;
#10 a = 42062; b = 53226; cin = 0;
#10 a = 55059; b = 4668; cin = 0;
#10 a = 15872; b = 13981; cin = 0;
#10 a = 55138; b = 39559; cin = 1;
#10 a = 6425; b = 51926; cin = 1;
#10 a = 6261; b = 57555; cin = 0;
#10 a = 2543; b = 60210; cin = 1;
#10 a = 2553; b = 26917; cin = 1;
#10 a = 46851; b = 67144; cin = 0;
#10 a = 40379; b = 38352; cin = 1;
#10 a = 5528; b = 56766; cin = 1;
#10 a = 42447; b = 41826; cin = 1;
#10 a = 8931; b = 34050; cin = 0;
#10 a = 40844; b = 19189; cin = 1;
#10 a = 38577; b = 1966; cin = 1;
#10 a = 46192; b = 8227; cin = 0;
#10 a = 52906; b = 57123; cin = 1;
#10 a = 31256; b = 59676; cin = 0;
#10 a = 41015; b = 36527; cin = 0;
#10 a = 54185; b = 53259; cin = 1;
#10 a = 3296; b = 58787; cin = 1;
#10 a = 5633; b = 7586; cin = 1;
#10 a = 58991; b = 62870; cin = 0;
#10 a = 32681; b = 33714; cin = 1;
#10 a = 45931; b = 48643; cin = 1;
#10 a = 17458; b = 1188; cin = 1;
#10 a = 46541; b = 54094; cin = 0;
#10 a = 42186; b = 61702; cin = 0;
#10 a = 64748; b = 32717; cin = 0;
#10 a = 60807; b = 16902; cin = 1;
#10 a = 1570; b = 20198; cin = 0;
#10 a = 45451; b = 2184; cin = 1;
#10 a = 14807; b = 37527; cin = 1;
#10 a = 64565; b = 208; cin = 1;
#10 a = 63512; b = 22491; cin = 0;
#10 a = 64425; b = 39950; cin = 0;
#10 a = 49918; b = 62843; cin = 1;
#10 a = 22534; b = 35029; cin = 1;
#10 a = 31179; b = 6129; cin = 1;
#10 a = 6351; b = 43288; cin = 1;
#10 a = 57486; b = 44858; cin = 0;
#10 a = 27408; b = 66662; cin = 0;
#10 a = 51269; b = 11469; cin = 1;
#10 a = 68000; b = 6034; cin = 1;
#10 a = 24797; b = 45898; cin = 1;
#10 a = 30238; b = 40323; cin = 1;
#10 a = 60514; b = 66594; cin = 0;
#10 a = 51237; b = 19128; cin = 1;
#10 a = 33663; b = 50307; cin = 0;
#10 a = 48806; b = 33010; cin = 1;
#10 a = 33555; b = 66848; cin = 1;
#10 a = 38503; b = 609; cin = 1;
#10 a = 45635; b = 51878; cin = 0;
#10 a = 66646; b = 26231; cin = 0;
#10 a = 64218; b = 27380; cin = 0;
#10 a = 14281; b = 57618; cin = 0;
#10 a = 50646; b = 24485; cin = 0;
#10 a = 56206; b = 5722; cin = 0;
#10 a = 50443; b = 39385; cin = 0;
#10 a = 27161; b = 64543; cin = 0;
#10 a = 47168; b = 28099; cin = 1;
#10 a = 18386; b = 42954; cin = 0;
#10 a = 56265; b = 64942; cin = 0;
#10 a = 11966; b = 37940; cin = 1;
#10 a = 20052; b = 32158; cin = 0;
#10 a = 4037; b = 22791; cin = 0;
#10 a = 28345; b = 49789; cin = 1;
#10 a = 25599; b = 35995; cin = 0;
#10 a = 41981; b = 62790; cin = 1;
#10 a = 15023; b = 66304; cin = 1;
#10 a = 67428; b = 19824; cin = 0;
#10 a = 23033; b = 14562; cin = 0;
#10 a = 2895; b = 828; cin = 0;
#10 a = 57339; b = 59146; cin = 1;
#10 a = 68015; b = 9198; cin = 1;
#10 a = 36071; b = 13235; cin = 1;
#10 a = 38097; b = 17932; cin = 0;
#10 a = 64609; b = 43531; cin = 0;
#10 a = 26843; b = 61865; cin = 0;
#10 a = 51166; b = 53240; cin = 0;
#10 a = 33; b = 27020; cin = 1;
#10 a = 46999; b = 50053; cin = 1;
#10 a = 43272; b = 29300; cin = 1;
#10 a = 34486; b = 16640; cin = 1;
#10 a = 63641; b = 14655; cin = 0;
#10 a = 31307; b = 27078; cin = 1;
#10 a = 21764; b = 65175; cin = 0;
#10 a = 38362; b = 36136; cin = 1;
#10 a = 67308; b = 39331; cin = 0;
#10 a = 65397; b = 20498; cin = 1;
#10 a = 59789; b = 20531; cin = 1;
#10 a = 50358; b = 43883; cin = 1;
#10 a = 9138; b = 63507; cin = 1;
#10 a = 61449; b = 27993; cin = 1;
#10 a = 32907; b = 67987; cin = 0;
#10 a = 13563; b = 29294; cin = 0;
#10 a = 53806; b = 27410; cin = 0;
#10 a = 18334; b = 42124; cin = 0;
#10 a = 26394; b = 15785; cin = 0;
#10 a = 2670; b = 11182; cin = 0;
#10 a = 32187; b = 47323; cin = 1;
#10 a = 18725; b = 27682; cin = 0;
#10 a = 55316; b = 13172; cin = 1;
#10 a = 51207; b = 4621; cin = 1;
#10 a = 40091; b = 37528; cin = 0;
#10 a = 43629; b = 27443; cin = 0;
#10 a = 4246; b = 57602; cin = 0;
#10 a = 52742; b = 5936; cin = 0;
#10 a = 21022; b = 32330; cin = 1;
#10 a = 4986; b = 11353; cin = 1;
#10 a = 55800; b = 43540; cin = 1;
#10 a = 57146; b = 62265; cin = 1;
#10 a = 32374; b = 47581; cin = 1;
#10 a = 47462; b = 5141; cin = 0;
#10 a = 20543; b = 45232; cin = 1;
#10 a = 37963; b = 65213; cin = 0;
#10 a = 14677; b = 69459; cin = 0;
#10 a = 18801; b = 52201; cin = 1;
#10 a = 41401; b = 49576; cin = 1;
#10 a = 56139; b = 30914; cin = 0;
#10 a = 35706; b = 63067; cin = 1;
#10 a = 38949; b = 50213; cin = 0;
#10 a = 46226; b = 58939; cin = 0;
#10 a = 66675; b = 36401; cin = 1;
#10 a = 21746; b = 33296; cin = 1;
#10 a = 37049; b = 1259; cin = 0;
#10 a = 9795; b = 15936; cin = 0;
#10 a = 16496; b = 11089; cin = 1;
#10 a = 52781; b = 28843; cin = 1;
#10 a = 4100; b = 14982; cin = 0;
#10 a = 36773; b = 27040; cin = 1;
#10 a = 19338; b = 65990; cin = 0;
#10 a = 64168; b = 42216; cin = 1;
#10 a = 62932; b = 38892; cin = 1;
#10 a = 43189; b = 36990; cin = 1;
#10 a = 68678; b = 50391; cin = 1;
#10 a = 19381; b = 36538; cin = 1;
#10 a = 15895; b = 53034; cin = 1;
#10 a = 40962; b = 12167; cin = 0;
#10 a = 21958; b = 16268; cin = 0;
#10 a = 33868; b = 29393; cin = 0;
#10 a = 15197; b = 48731; cin = 0;
#10 a = 23091; b = 42899; cin = 1;
#10 a = 19924; b = 12184; cin = 1;
#10 a = 29511; b = 55373; cin = 1;
#10 a = 2395; b = 54052; cin = 0;
#10 a = 22890; b = 49785; cin = 0;
#10 a = 35673; b = 42032; cin = 1;
#10 a = 35898; b = 12994; cin = 0;
#10 a = 64966; b = 34952; cin = 0;
#10 a = 15368; b = 45172; cin = 1;
#10 a = 62811; b = 36721; cin = 0;
#10 a = 36243; b = 59812; cin = 0;
#10 a = 4596; b = 9737; cin = 0;
#10 a = 58193; b = 15600; cin = 1;
#10 a = 8780; b = 64347; cin = 1;
#10 a = 56110; b = 17237; cin = 0;
#10 a = 46331; b = 29263; cin = 0;
#10 a = 43234; b = 41513; cin = 1;
#10 a = 28656; b = 36480; cin = 1;
#10 a = 6699; b = 51848; cin = 0;
#10 a = 14134; b = 44659; cin = 1;
#10 a = 46653; b = 57255; cin = 0;
#10 a = 28423; b = 38203; cin = 1;
#10 a = 22377; b = 26397; cin = 1;
#10 a = 1704; b = 11529; cin = 1;
#10 a = 11436; b = 43992; cin = 0;
#10 a = 47304; b = 20323; cin = 1;
#10 a = 55205; b = 39909; cin = 1;
#10 a = 6100; b = 68565; cin = 1;
#10 a = 14651; b = 51616; cin = 1;
#10 a = 68375; b = 42103; cin = 1;
#10 a = 65173; b = 18756; cin = 0;
#10 a = 51783; b = 47179; cin = 1;
#10 a = 834; b = 69556; cin = 0;
#10 a = 35485; b = 47612; cin = 0;
#10 a = 18132; b = 35400; cin = 0;
#10 a = 40721; b = 12705; cin = 1;
#10 a = 68924; b = 44262; cin = 0;
#10 a = 22289; b = 50362; cin = 1;
#10 a = 34838; b = 41365; cin = 0;
#10 a = 52884; b = 39741; cin = 1;
#10 a = 68293; b = 11266; cin = 1;
#10 a = 957; b = 39401; cin = 0;
#10 a = 18176; b = 40235; cin = 0;
#10 a = 61793; b = 5720; cin = 0;
#10 a = 23291; b = 205; cin = 1;
#10 a = 28781; b = 17278; cin = 0;
#10 a = 30946; b = 16202; cin = 0;
#10 a = 3020; b = 14844; cin = 0;
#10 a = 20011; b = 49682; cin = 1;
#10 a = 18619; b = 8918; cin = 0;
#10 a = 35682; b = 53563; cin = 0;
#10 a = 1501; b = 30872; cin = 1;
#10 a = 14499; b = 49049; cin = 0;
#10 a = 3405; b = 17194; cin = 1;
#10 a = 39924; b = 40485; cin = 0;
#10 a = 41843; b = 69266; cin = 0;
#10 a = 32819; b = 30212; cin = 0;
#10 a = 68057; b = 33232; cin = 0;
#10 a = 60009; b = 53243; cin = 1;
#10 a = 23326; b = 48215; cin = 1;
#10 a = 26385; b = 13897; cin = 1;
#10 a = 17061; b = 15399; cin = 1;
#10 a = 47139; b = 6250; cin = 0;
#10 a = 23803; b = 56008; cin = 0;
#10 a = 52540; b = 25932; cin = 1;
#10 a = 57834; b = 44127; cin = 1;
#10 a = 10406; b = 53298; cin = 1;
#10 a = 25533; b = 51355; cin = 1;
#10 a = 31855; b = 41364; cin = 1;
#10 a = 64212; b = 64690; cin = 0;
#10 a = 35488; b = 67427; cin = 1;
#10 a = 60327; b = 60841; cin = 0;
#10 a = 22390; b = 14332; cin = 1;
#10 a = 33503; b = 38135; cin = 1;
#10 a = 38161; b = 67028; cin = 1;
#10 a = 36953; b = 54862; cin = 0;
#10 a = 57714; b = 41621; cin = 0;
#10 a = 38688; b = 67154; cin = 1;
#10 a = 52893; b = 5361; cin = 1;
#10 a = 3046; b = 69574; cin = 1;
#10 a = 1414; b = 35062; cin = 1;
#10 a = 60032; b = 1741; cin = 0;
#10 a = 64048; b = 24131; cin = 0;
#10 a = 27019; b = 33986; cin = 1;
#10 a = 69646; b = 2148; cin = 1;
#10 a = 44557; b = 15453; cin = 0;
#10 a = 39947; b = 3167; cin = 1;
#10 a = 18635; b = 41855; cin = 1;
#10 a = 25030; b = 1101; cin = 0;
#10 a = 2789; b = 50499; cin = 0;
#10 a = 67943; b = 51914; cin = 0;
#10 a = 36876; b = 18298; cin = 1;
#10 a = 66650; b = 58698; cin = 1;
#10 a = 40756; b = 15718; cin = 1;
#10 a = 29349; b = 15364; cin = 1;
#10 a = 14971; b = 59922; cin = 0;
#10 a = 31807; b = 29869; cin = 0;
#10 a = 20264; b = 48505; cin = 1;
#10 a = 52227; b = 3535; cin = 0;
#10 a = 65903; b = 52677; cin = 0;
#10 a = 9154; b = 26972; cin = 0;
#10 a = 33818; b = 63848; cin = 0;
#10 a = 36576; b = 60498; cin = 0;
#10 a = 63465; b = 7606; cin = 0;
#10 a = 54340; b = 36955; cin = 1;
#10 a = 23716; b = 51926; cin = 1;
#10 a = 8544; b = 60085; cin = 0;
#10 a = 66540; b = 10349; cin = 1;
#10 a = 26392; b = 38928; cin = 1;
#10 a = 33696; b = 34832; cin = 0;
#10 a = 21500; b = 43986; cin = 0;
#10 a = 37570; b = 7804; cin = 0;
#10 a = 25586; b = 20732; cin = 0;
#10 a = 48653; b = 14197; cin = 0;
#10 a = 17437; b = 44890; cin = 1;
#10 a = 1586; b = 44958; cin = 0;
#10 a = 22009; b = 53502; cin = 1;
#10 a = 48654; b = 50043; cin = 1;
#10 a = 53803; b = 52787; cin = 1;
#10 a = 38840; b = 62835; cin = 1;
#10 a = 52906; b = 14336; cin = 1;
#10 a = 23944; b = 28258; cin = 0;
#10 a = 35182; b = 30197; cin = 0;
#10 a = 13270; b = 8850; cin = 0;
#10 a = 68964; b = 2639; cin = 0;
#10 a = 21614; b = 50578; cin = 0;
#10 a = 2542; b = 2587; cin = 0;
#10 a = 19907; b = 51241; cin = 1;
#10 a = 47622; b = 35045; cin = 0;
#10 a = 44266; b = 50237; cin = 0;
#10 a = 5741; b = 33144; cin = 0;
#10 a = 11203; b = 33440; cin = 0;
#10 a = 821; b = 44975; cin = 1;
#10 a = 57523; b = 58245; cin = 1;
#10 a = 58423; b = 33562; cin = 1;
#10 a = 34213; b = 55176; cin = 1;
#10 a = 31313; b = 34070; cin = 0;
#10 a = 11916; b = 53977; cin = 0;
#10 a = 65265; b = 31600; cin = 1;
#10 a = 55050; b = 5866; cin = 0;
#10 a = 14022; b = 57959; cin = 0;
#10 a = 33682; b = 69162; cin = 1;
#10 a = 57952; b = 46335; cin = 0;
#10 a = 66068; b = 33859; cin = 1;
#10 a = 59385; b = 22282; cin = 1;
#10 a = 31694; b = 32848; cin = 1;
#10 a = 54581; b = 40513; cin = 1;
#10 a = 10056; b = 28781; cin = 1;
#10 a = 63124; b = 24047; cin = 1;
#10 a = 57589; b = 55449; cin = 1;
#10 a = 32291; b = 45823; cin = 0;
#10 a = 16490; b = 55857; cin = 1;
#10 a = 10481; b = 43809; cin = 0;
#10 a = 49447; b = 16229; cin = 1;
#10 a = 6658; b = 5615; cin = 0;
#10 a = 43784; b = 13661; cin = 0;
#10 a = 42437; b = 68243; cin = 1;
#10 a = 5161; b = 8299; cin = 1;
#10 a = 68214; b = 47775; cin = 0;
#10 a = 69219; b = 35364; cin = 1;
#10 a = 52442; b = 44007; cin = 0;
#10 a = 69976; b = 60497; cin = 1;
#10 a = 40321; b = 47330; cin = 0;
#10 a = 9706; b = 26777; cin = 0;
#10 a = 36597; b = 33436; cin = 1;
#10 a = 38475; b = 53572; cin = 0;
#10 a = 3201; b = 26009; cin = 1;
#10 a = 31145; b = 31170; cin = 0;
#10 a = 41518; b = 5736; cin = 1;
#10 a = 28642; b = 51307; cin = 1;
#10 a = 1215; b = 10101; cin = 1;
#10 a = 19611; b = 10078; cin = 0;
#10 a = 23864; b = 26751; cin = 1;
#10 a = 48278; b = 36457; cin = 0;
#10 a = 18922; b = 49407; cin = 0;
#10 a = 41533; b = 17882; cin = 0;
#10 a = 7806; b = 67436; cin = 0;
#10 a = 42321; b = 28581; cin = 0;
#10 a = 61488; b = 46451; cin = 1;
#10 a = 34781; b = 5093; cin = 0;
#10 a = 43439; b = 6308; cin = 0;
#10 a = 26104; b = 2271; cin = 0;
#10 a = 21970; b = 26135; cin = 1;
#10 a = 18815; b = 50765; cin = 1;
#10 a = 42438; b = 69688; cin = 0;
#10 a = 5848; b = 41221; cin = 0;
#10 a = 69183; b = 25379; cin = 0;
#10 a = 42175; b = 67701; cin = 1;
#10 a = 69041; b = 35541; cin = 0;
#10 a = 31644; b = 46674; cin = 1;
#10 a = 45555; b = 20113; cin = 1;
#10 a = 45919; b = 22569; cin = 0;
#10 a = 56361; b = 44540; cin = 1;
#10 a = 69906; b = 39707; cin = 1;
#10 a = 26261; b = 12145; cin = 1;
#10 a = 32023; b = 64346; cin = 0;
#10 a = 32020; b = 63529; cin = 0;
#10 a = 5804; b = 12056; cin = 1;
#10 a = 8170; b = 11097; cin = 0;
#10 a = 9690; b = 42742; cin = 0;
#10 a = 16304; b = 64649; cin = 0;
#10 a = 5577; b = 40568; cin = 1;
#10 a = 43474; b = 3281; cin = 1;
#10 a = 37505; b = 3187; cin = 1;
#10 a = 58654; b = 5801; cin = 0;
#10 a = 9491; b = 37824; cin = 0;
#10 a = 47902; b = 69844; cin = 1;
#10 a = 18044; b = 5649; cin = 1;
#10 a = 55887; b = 60171; cin = 1;
#10 a = 35623; b = 69861; cin = 1;
#10 a = 62033; b = 62517; cin = 0;
#10 a = 14909; b = 44447; cin = 0;
#10 a = 60355; b = 17921; cin = 1;
#10 a = 33044; b = 31778; cin = 0;
#10 a = 69089; b = 20433; cin = 1;
#10 a = 23632; b = 6276; cin = 0;
#10 a = 18872; b = 30530; cin = 0;
#10 a = 53994; b = 48574; cin = 1;
#10 a = 31171; b = 10813; cin = 0;
#10 a = 65798; b = 46436; cin = 0;
#10 a = 49519; b = 14822; cin = 1;
#10 a = 27889; b = 29731; cin = 0;
#10 a = 46827; b = 66438; cin = 1;
#10 a = 45398; b = 5835; cin = 0;
#10 a = 23509; b = 4924; cin = 1;
#10 a = 53772; b = 4908; cin = 1;
#10 a = 5508; b = 133; cin = 0;
#10 a = 3441; b = 54127; cin = 0;
#10 a = 53374; b = 61650; cin = 0;
#10 a = 69831; b = 57449; cin = 0;
#10 a = 16149; b = 36968; cin = 0;
#10 a = 1336; b = 64858; cin = 0;
#10 a = 30971; b = 18037; cin = 0;
#10 a = 31230; b = 39788; cin = 1;
#10 a = 63268; b = 39649; cin = 0;
#10 a = 22091; b = 23421; cin = 0;
#10 a = 57191; b = 5282; cin = 1;
#10 a = 52821; b = 55075; cin = 0;
#10 a = 3377; b = 38449; cin = 1;
#10 a = 34747; b = 38280; cin = 0;
#10 a = 18906; b = 30781; cin = 0;
#10 a = 17886; b = 32118; cin = 0;
#10 a = 22950; b = 39441; cin = 0;
#10 a = 24453; b = 671; cin = 0;
#10 a = 8142; b = 63940; cin = 1;
#10 a = 43108; b = 16031; cin = 0;
#10 a = 12983; b = 3222; cin = 0;
#10 a = 52990; b = 32395; cin = 1;
#10 a = 29829; b = 35773; cin = 1;
#10 a = 68318; b = 520; cin = 1;
#10 a = 608; b = 19426; cin = 1;
#10 a = 16218; b = 37313; cin = 1;
#10 a = 3039; b = 36615; cin = 0;
#10 a = 7897; b = 61068; cin = 1;
#10 a = 28895; b = 45563; cin = 1;
#10 a = 65894; b = 18671; cin = 1;
#10 a = 56314; b = 31654; cin = 1;
#10 a = 28369; b = 60997; cin = 1;
#10 a = 55498; b = 67178; cin = 0;
#10 a = 27429; b = 65496; cin = 0;
#10 a = 13993; b = 42456; cin = 1;
#10 a = 31338; b = 58674; cin = 0;
#10 a = 57153; b = 61713; cin = 1;
#10 a = 52409; b = 45962; cin = 0;
#10 a = 24688; b = 4857; cin = 1;
#10 a = 37260; b = 751; cin = 0;
#10 a = 65863; b = 33418; cin = 1;
#10 a = 50392; b = 38139; cin = 0;
#10 a = 20965; b = 23637; cin = 0;
#10 a = 3663; b = 27419; cin = 0;
#10 a = 33234; b = 41412; cin = 0;
#10 a = 12231; b = 49102; cin = 0;
#10 a = 4893; b = 12607; cin = 0;
#10 a = 34170; b = 65016; cin = 0;
#10 a = 30868; b = 66056; cin = 0;
#10 a = 49481; b = 33316; cin = 1;
#10 a = 16766; b = 5531; cin = 1;
#10 a = 62057; b = 55924; cin = 0;
#10 a = 28345; b = 53241; cin = 0;
#10 a = 14515; b = 33257; cin = 1;
#10 a = 19829; b = 42843; cin = 1;
#10 a = 20303; b = 55074; cin = 1;
#10 a = 9451; b = 36319; cin = 0;
#10 a = 13017; b = 46841; cin = 0;
#10 a = 16194; b = 7710; cin = 0;
#10 a = 580; b = 57191; cin = 1;
#10 a = 8421; b = 3957; cin = 0;
#10 a = 49681; b = 42366; cin = 0;
#10 a = 59079; b = 47063; cin = 0;
#10 a = 68467; b = 61578; cin = 1;
#10 a = 35274; b = 57759; cin = 0;
#10 a = 19845; b = 8062; cin = 0;
#10 a = 53518; b = 63866; cin = 1;
#10 a = 29798; b = 6883; cin = 0;
#10 a = 47446; b = 69429; cin = 0;
#10 a = 61151; b = 46361; cin = 0;
#10 a = 60876; b = 54783; cin = 1;
#10 a = 66132; b = 34464; cin = 0;
#10 a = 57313; b = 23543; cin = 1;
#10 a = 54439; b = 22011; cin = 0;
#10 a = 61174; b = 33637; cin = 1;
#10 a = 40752; b = 53483; cin = 0;
#10 a = 5404; b = 37001; cin = 0;
#10 a = 29079; b = 66800; cin = 1;
#10 a = 53243; b = 20598; cin = 1;
#10 a = 61470; b = 58101; cin = 0;
#10 a = 33240; b = 48977; cin = 1;
#10 a = 8967; b = 45110; cin = 1;
#10 a = 3413; b = 8775; cin = 1;
#10 a = 44923; b = 39566; cin = 0;
#10 a = 31659; b = 30740; cin = 1;
#10 a = 52506; b = 1492; cin = 0;
#10 a = 57768; b = 53248; cin = 0;
#10 a = 56896; b = 12327; cin = 0;
#10 a = 62908; b = 41922; cin = 0;
#10 a = 68349; b = 33392; cin = 0;
#10 a = 26503; b = 42984; cin = 1;
#10 a = 63089; b = 28304; cin = 1;
#10 a = 16842; b = 31717; cin = 0;
#10 a = 17787; b = 6640; cin = 0;
#10 a = 63447; b = 14651; cin = 0;
#10 a = 2745; b = 43510; cin = 0;
#10 a = 41877; b = 31278; cin = 0;
#10 a = 1659; b = 18175; cin = 1;
#10 a = 50945; b = 11083; cin = 0;
#10 a = 50830; b = 55784; cin = 0;
#10 a = 38816; b = 12287; cin = 1;
#10 a = 52131; b = 51728; cin = 1;
#10 a = 40557; b = 68571; cin = 0;
#10 a = 60461; b = 62710; cin = 1;
#10 a = 3580; b = 32510; cin = 0;
#10 a = 142; b = 35255; cin = 0;
#10 a = 68197; b = 53484; cin = 1;
#10 a = 49499; b = 55144; cin = 0;
#10 a = 19481; b = 12441; cin = 1;
#10 a = 31385; b = 63271; cin = 1;
#10 a = 53033; b = 32087; cin = 0;
#10 a = 24018; b = 60571; cin = 1;
#10 a = 23307; b = 31128; cin = 0;
#10 a = 54314; b = 67941; cin = 0;
#10 a = 68313; b = 1521; cin = 0;
#10 a = 26963; b = 48016; cin = 1;
#10 a = 29124; b = 46213; cin = 0;
#10 a = 38915; b = 25712; cin = 0;
#10 a = 20529; b = 45193; cin = 1;
#10 a = 35930; b = 52930; cin = 1;
#10 a = 37115; b = 12316; cin = 0;
#10 a = 50587; b = 36334; cin = 1;
#10 a = 22140; b = 59642; cin = 1;
#10 a = 62264; b = 20308; cin = 1;
#10 a = 1451; b = 18621; cin = 0;
#10 a = 19499; b = 45584; cin = 0;
#10 a = 2803; b = 51060; cin = 1;
#10 a = 39591; b = 19975; cin = 0;
#10 a = 37875; b = 16856; cin = 1;
#10 a = 48600; b = 52786; cin = 0;
#10 a = 28949; b = 19901; cin = 0;
#10 a = 41386; b = 489; cin = 0;
#10 a = 44393; b = 68981; cin = 0;
#10 a = 31233; b = 37598; cin = 0;
#10 a = 39662; b = 15401; cin = 1;
#10 a = 25964; b = 34900; cin = 0;
#10 a = 60283; b = 37703; cin = 0;
#10 a = 47166; b = 53646; cin = 0;
#10 a = 59762; b = 21521; cin = 0;
#10 a = 23904; b = 46474; cin = 1;
#10 a = 40976; b = 5423; cin = 0;
#10 a = 46716; b = 23161; cin = 1;
#10 a = 18790; b = 43907; cin = 1;
#10 a = 3211; b = 5140; cin = 1;
#10 a = 31587; b = 21154; cin = 0;
#10 a = 54937; b = 47118; cin = 0;
#10 a = 30223; b = 13753; cin = 0;
#10 a = 32921; b = 60920; cin = 0;
#10 a = 9243; b = 27034; cin = 0;
#10 a = 2422; b = 50938; cin = 0;
#10 a = 24739; b = 21914; cin = 1;
#10 a = 66957; b = 68630; cin = 1;
#10 a = 16017; b = 63773; cin = 0;
#10 a = 34058; b = 66984; cin = 0;
#10 a = 66049; b = 4923; cin = 0;
#10 a = 67089; b = 36212; cin = 0;
#10 a = 9381; b = 42787; cin = 0;
#10 a = 35729; b = 5709; cin = 0;
#10 a = 45724; b = 14952; cin = 0;
#10 a = 7240; b = 63726; cin = 1;
#10 a = 61582; b = 64817; cin = 1;
#10 a = 27699; b = 38127; cin = 0;
#10 a = 63330; b = 54144; cin = 1;
#10 a = 2868; b = 64554; cin = 1;
#10 a = 17546; b = 60603; cin = 0;
#10 a = 53378; b = 57692; cin = 1;
#10 a = 19033; b = 43425; cin = 0;
#10 a = 22089; b = 9155; cin = 1;
#10 a = 38769; b = 54879; cin = 0;
#10 a = 12483; b = 38471; cin = 0;
#10 a = 37136; b = 6405; cin = 0;
#10 a = 60056; b = 10456; cin = 1;
#10 a = 57958; b = 3787; cin = 1;
#10 a = 49633; b = 6655; cin = 1;
#10 a = 14644; b = 24202; cin = 0;
#10 a = 30930; b = 53932; cin = 0;
#10 a = 13429; b = 2965; cin = 1;
#10 a = 38716; b = 1406; cin = 0;
#10 a = 69711; b = 40175; cin = 1;
#10 a = 68363; b = 29011; cin = 0;
#10 a = 60742; b = 66147; cin = 1;
#10 a = 47938; b = 56203; cin = 0;
#10 a = 3261; b = 44161; cin = 1;
#10 a = 59080; b = 146; cin = 0;
#10 a = 15805; b = 61142; cin = 0;
#10 a = 56781; b = 22073; cin = 1;
#10 a = 38153; b = 35502; cin = 0;
#10 a = 62950; b = 4218; cin = 1;
#10 a = 3255; b = 50282; cin = 0;
#10 a = 44790; b = 48645; cin = 1;
#10 a = 54797; b = 15739; cin = 1;
#10 a = 1208; b = 63677; cin = 0;
#10 a = 28076; b = 43290; cin = 0;
#10 a = 35083; b = 8722; cin = 0;
#10 a = 48746; b = 24527; cin = 1;
#10 a = 16610; b = 57660; cin = 0;
#10 a = 61111; b = 2165; cin = 0;
#10 a = 38578; b = 41468; cin = 1;
#10 a = 63803; b = 21075; cin = 1;
#10 a = 59203; b = 65865; cin = 0;
#10 a = 59967; b = 50662; cin = 0;
#10 a = 56878; b = 28223; cin = 1;
#10 a = 39992; b = 32651; cin = 0;
#10 a = 19972; b = 67735; cin = 0;
#10 a = 99; b = 46481; cin = 0;
#10 a = 41368; b = 39443; cin = 0;
#10 a = 34710; b = 30555; cin = 0;
#10 a = 39906; b = 69133; cin = 0;
#10 a = 25673; b = 39288; cin = 1;
#10 a = 61722; b = 28491; cin = 0;
#10 a = 52769; b = 64810; cin = 1;
#10 a = 35907; b = 51688; cin = 0;
#10 a = 36370; b = 68033; cin = 1;
#10 a = 32828; b = 18005; cin = 0;
#10 a = 61657; b = 18104; cin = 1;
#10 a = 21365; b = 59472; cin = 1;
#10 a = 15085; b = 534; cin = 0;
#10 a = 34619; b = 40441; cin = 1;
#10 a = 1973; b = 66114; cin = 1;
#10 a = 60402; b = 34189; cin = 0;
#10 a = 44697; b = 63310; cin = 1;
#10 a = 32358; b = 29217; cin = 1;
#10 a = 48242; b = 41939; cin = 0;
#10 a = 26777; b = 4768; cin = 0;
#10 a = 49400; b = 66425; cin = 0;
#10 a = 48503; b = 64142; cin = 1;
#10 a = 63402; b = 9227; cin = 1;
#10 a = 38856; b = 20199; cin = 0;
#10 a = 59795; b = 22172; cin = 1;
#10 a = 50022; b = 58927; cin = 0;
#10 a = 45093; b = 9976; cin = 0;
#10 a = 34974; b = 42334; cin = 1;
#10 a = 52895; b = 66928; cin = 0;
#10 a = 22498; b = 23705; cin = 0;
#10 a = 56458; b = 3105; cin = 1;
#10 a = 38522; b = 27961; cin = 1;
#10 a = 56411; b = 21363; cin = 1;
#10 a = 28483; b = 60220; cin = 0;
#10 a = 63699; b = 50015; cin = 0;
#10 a = 48678; b = 6390; cin = 1;
#10 a = 44198; b = 27835; cin = 1;
#10 a = 33028; b = 39161; cin = 1;
#10 a = 27427; b = 22056; cin = 1;
#10 a = 17414; b = 20906; cin = 1;
#10 a = 12168; b = 7364; cin = 0;
#10 a = 26052; b = 22239; cin = 1;
#10 a = 34077; b = 8650; cin = 1;
#10 a = 51330; b = 13485; cin = 1;
#10 a = 65134; b = 7185; cin = 0;
#10 a = 31111; b = 32215; cin = 0;
#10 a = 8718; b = 52766; cin = 1;
#10 a = 19950; b = 62146; cin = 0;
#10 a = 49867; b = 19574; cin = 1;
#10 a = 53065; b = 36988; cin = 1;
#10 a = 33616; b = 25508; cin = 0;
#10 a = 39976; b = 27912; cin = 1;
#10 a = 27946; b = 61990; cin = 1;
#10 a = 13631; b = 43320; cin = 1;
#10 a = 59536; b = 14807; cin = 0;
#10 a = 61808; b = 45918; cin = 1;
#10 a = 46823; b = 54636; cin = 1;
#10 a = 13320; b = 50938; cin = 0;
#10 a = 65331; b = 7158; cin = 0;
#10 a = 45750; b = 60223; cin = 0;
#10 a = 47075; b = 191; cin = 0;
#10 a = 55765; b = 40167; cin = 1;
#10 a = 63046; b = 44465; cin = 1;
#10 a = 31682; b = 58096; cin = 1;
#10 a = 13803; b = 23984; cin = 0;
#10 a = 49461; b = 15793; cin = 0;
#10 a = 23686; b = 62616; cin = 1;
#10 a = 50678; b = 52288; cin = 1;
#10 a = 46168; b = 23971; cin = 1;
#10 a = 37584; b = 69721; cin = 0;
#10 a = 42340; b = 46797; cin = 1;
#10 a = 48956; b = 8914; cin = 1;
#10 a = 37133; b = 48313; cin = 0;
#10 a = 63652; b = 9995; cin = 1;
#10 a = 39844; b = 23798; cin = 1;
#10 a = 30842; b = 3259; cin = 0;
#10 a = 44111; b = 26945; cin = 0;
#10 a = 18368; b = 53975; cin = 1;
#10 a = 19915; b = 6495; cin = 0;
#10 a = 28621; b = 44079; cin = 0;
#10 a = 27549; b = 62771; cin = 1;
#10 a = 3021; b = 41728; cin = 1;
#10 a = 18660; b = 55213; cin = 0;
#10 a = 55116; b = 25218; cin = 1;
#10 a = 9669; b = 65062; cin = 1;
#10 a = 58207; b = 2256; cin = 0;
#10 a = 28889; b = 22719; cin = 0;
#10 a = 38540; b = 17439; cin = 1;
#10 a = 30479; b = 37355; cin = 1;
#10 a = 46389; b = 65976; cin = 0;
#10 a = 38373; b = 69877; cin = 0;
#10 a = 53506; b = 2898; cin = 0;
#10 a = 53906; b = 67910; cin = 1;
#10 a = 32618; b = 53027; cin = 1;
#10 a = 21326; b = 62696; cin = 1;
#10 a = 56535; b = 27255; cin = 0;
#10 a = 25004; b = 56145; cin = 1;
#10 a = 66770; b = 24685; cin = 1;
#10 a = 68863; b = 55164; cin = 0;
#10 a = 7452; b = 7905; cin = 0;
#10 a = 36473; b = 46279; cin = 1;
#10 a = 58265; b = 6137; cin = 0;
#10 a = 51785; b = 60043; cin = 0;
#10 a = 6870; b = 22662; cin = 1;
#10 a = 57174; b = 20340; cin = 0;
#10 a = 32539; b = 6875; cin = 1;
#10 a = 32865; b = 31879; cin = 0;
#10 a = 9559; b = 5001; cin = 1;
#10 a = 26396; b = 3865; cin = 1;
#10 a = 34236; b = 11317; cin = 1;
#10 a = 60756; b = 47790; cin = 0;
#10 a = 17153; b = 12407; cin = 1;
#10 a = 22801; b = 40544; cin = 1;
#10 a = 2712; b = 47415; cin = 1;
#10 a = 59297; b = 34589; cin = 1;
#10 a = 14931; b = 43480; cin = 0;
#10 a = 67821; b = 52698; cin = 0;
#10 a = 13207; b = 62257; cin = 1;
#10 a = 29631; b = 18653; cin = 0;
#10 a = 31218; b = 29241; cin = 0;
#10 a = 40711; b = 66349; cin = 0;
#10 a = 26483; b = 59854; cin = 0;
#10 a = 64745; b = 59008; cin = 0;
#10 a = 23050; b = 61720; cin = 1;
#10 a = 4017; b = 51017; cin = 0;
#10 a = 5324; b = 42301; cin = 1;
#10 a = 13506; b = 16474; cin = 1;
#10 a = 29920; b = 6033; cin = 0;
#10 a = 51336; b = 35664; cin = 1;
#10 a = 6616; b = 66883; cin = 0;
#10 a = 19566; b = 37594; cin = 1;
#10 a = 10307; b = 40430; cin = 1;
#10 a = 59807; b = 35175; cin = 1;
#10 a = 9851; b = 58225; cin = 1;
#10 a = 7311; b = 62242; cin = 1;
#10 a = 15711; b = 43918; cin = 0;
#10 a = 43944; b = 57424; cin = 0;
#10 a = 54875; b = 17345; cin = 1;
#10 a = 10767; b = 68681; cin = 0;
#10 a = 55312; b = 51649; cin = 1;
#10 a = 59098; b = 1216; cin = 1;
#10 a = 35585; b = 57875; cin = 1;
#10 a = 1927; b = 24034; cin = 0;
#10 a = 3628; b = 33885; cin = 1;
#10 a = 20698; b = 41196; cin = 1;
#10 a = 65137; b = 33260; cin = 1;
#10 a = 58229; b = 53556; cin = 0;
#10 a = 44147; b = 14784; cin = 1;
#10 a = 12450; b = 25551; cin = 0;
#10 a = 16418; b = 10864; cin = 1;
#10 a = 63621; b = 46314; cin = 1;
#10 a = 8419; b = 58252; cin = 0;
#10 a = 39998; b = 60179; cin = 0;
#10 a = 13105; b = 40159; cin = 0;
#10 a = 20788; b = 60857; cin = 0;
#10 a = 67066; b = 32346; cin = 0;
#10 a = 17261; b = 66927; cin = 1;
#10 a = 24881; b = 17426; cin = 1;
#10 a = 26198; b = 29877; cin = 0;
#10 a = 2548; b = 46295; cin = 0;
#10 a = 30548; b = 39917; cin = 1;
#10 a = 36115; b = 24688; cin = 1;
#10 a = 29558; b = 41038; cin = 0;
#10 a = 47034; b = 30495; cin = 1;
#10 a = 4748; b = 51284; cin = 1;
#10 a = 3659; b = 24702; cin = 1;
#10 a = 58533; b = 41963; cin = 1;
#10 a = 50612; b = 66845; cin = 1;
#10 a = 33827; b = 69395; cin = 0;
#10 a = 18946; b = 1944; cin = 0;
#10 a = 14928; b = 32492; cin = 1;
#10 a = 57225; b = 68607; cin = 1;
#10 a = 17774; b = 4517; cin = 1;
#10 a = 61206; b = 51552; cin = 1;
#10 a = 28446; b = 32652; cin = 1;
#10 a = 56543; b = 12663; cin = 1;
#10 a = 69690; b = 1197; cin = 0;
#10 a = 33413; b = 28161; cin = 1;
#10 a = 60915; b = 61989; cin = 1;
#10 a = 48293; b = 57287; cin = 1;
#10 a = 58319; b = 2215; cin = 1;
#10 a = 14614; b = 35793; cin = 0;
#10 a = 65597; b = 29919; cin = 0;
#10 a = 63971; b = 21126; cin = 0;
#10 a = 69192; b = 49572; cin = 0;
#10 a = 55697; b = 12467; cin = 0;
#10 a = 66904; b = 12157; cin = 1;
#10 a = 26426; b = 45571; cin = 0;
#10 a = 52794; b = 36486; cin = 1;
#10 a = 8557; b = 14779; cin = 0;
#10 a = 12616; b = 49451; cin = 0;
#10 a = 49167; b = 64065; cin = 1;
#10 a = 60677; b = 59663; cin = 0;
#10 a = 30353; b = 29986; cin = 0;
#10 a = 4285; b = 29178; cin = 0;
#10 a = 10870; b = 61227; cin = 1;
#10 a = 53766; b = 58131; cin = 1;
#10 a = 4211; b = 60909; cin = 0;
#10 a = 52817; b = 43703; cin = 0;
#10 a = 69765; b = 28612; cin = 1;
#10 a = 3999; b = 17580; cin = 0;
#10 a = 56801; b = 66747; cin = 0;
#10 a = 51748; b = 57425; cin = 1;
#10 a = 30263; b = 64130; cin = 1;
#10 a = 29903; b = 44768; cin = 1;
#10 a = 55468; b = 55638; cin = 0;
#10 a = 69851; b = 15756; cin = 1;
#10 a = 50040; b = 66319; cin = 0;
#10 a = 28504; b = 49136; cin = 0;
#10 a = 43454; b = 25253; cin = 0;
#10 a = 49536; b = 5605; cin = 1;
#10 a = 35068; b = 38758; cin = 0;
#10 a = 14666; b = 20507; cin = 1;
#10 a = 6631; b = 50770; cin = 0;
#10 a = 28582; b = 57025; cin = 0;
#10 a = 56063; b = 18845; cin = 0;
#10 a = 4771; b = 18697; cin = 0;
#10 a = 57962; b = 45089; cin = 1;
#10 a = 32063; b = 3594; cin = 1;
#10 a = 2571; b = 47048; cin = 1;
#10 a = 1691; b = 26584; cin = 0;
#10 a = 18392; b = 38005; cin = 0;
#10 a = 8193; b = 29023; cin = 1;
#10 a = 31770; b = 35655; cin = 1;
#10 a = 49478; b = 64237; cin = 1;
#10 a = 18306; b = 50301; cin = 0;
#10 a = 19124; b = 55072; cin = 1;
#10 a = 35698; b = 19387; cin = 1;
#10 a = 48591; b = 27802; cin = 1;
#10 a = 16973; b = 30373; cin = 1;
#10 a = 10608; b = 32064; cin = 0;
#10 a = 32552; b = 26809; cin = 1;
#10 a = 46902; b = 35002; cin = 0;
#10 a = 34464; b = 66772; cin = 1;
#10 a = 2795; b = 22603; cin = 1;
#10 a = 4504; b = 17261; cin = 0;
#10 a = 1411; b = 36386; cin = 0;
#10 a = 63366; b = 2084; cin = 1;
#10 a = 30411; b = 27028; cin = 1;
#10 a = 47402; b = 44001; cin = 0;
#10 a = 17794; b = 30961; cin = 1;
#10 a = 14770; b = 63513; cin = 0;
#10 a = 26103; b = 16767; cin = 0;
#10 a = 42811; b = 51231; cin = 0;
#10 a = 48823; b = 54027; cin = 1;
#10 a = 1776; b = 34883; cin = 1;
#10 a = 5030; b = 36294; cin = 1;
#10 a = 39708; b = 29661; cin = 1;
#10 a = 23774; b = 36424; cin = 1;
#10 a = 35641; b = 13827; cin = 0;
#10 a = 54234; b = 7973; cin = 1;
#10 a = 11243; b = 22743; cin = 0;
#10 a = 18709; b = 25198; cin = 0;
#10 a = 13881; b = 68009; cin = 1;
#10 a = 29473; b = 23184; cin = 0;
#10 a = 20373; b = 1312; cin = 0;
#10 a = 52182; b = 6342; cin = 0;
#10 a = 26729; b = 46051; cin = 1;
#10 a = 26064; b = 46177; cin = 0;
#10 a = 6076; b = 11818; cin = 1;
#10 a = 6440; b = 42404; cin = 0;
#10 a = 37766; b = 53647; cin = 1;
#10 a = 62604; b = 48708; cin = 1;
#10 a = 34210; b = 62589; cin = 0;
#10 a = 33400; b = 68415; cin = 1;
#10 a = 16616; b = 18788; cin = 1;
#10 a = 34716; b = 970; cin = 0;
#10 a = 65463; b = 4051; cin = 1;
#10 a = 55870; b = 30115; cin = 0;
#10 a = 59054; b = 12543; cin = 0;
#10 a = 52417; b = 18984; cin = 1;
#10 a = 53753; b = 56750; cin = 0;
#10 a = 7832; b = 25706; cin = 1;
#10 a = 33461; b = 36269; cin = 0;
#10 a = 33452; b = 69669; cin = 1;
#10 a = 56627; b = 62637; cin = 1;
#10 a = 57466; b = 27354; cin = 1;
#10 a = 18296; b = 69169; cin = 0;
#10 a = 47881; b = 55039; cin = 0;
#10 a = 7291; b = 20446; cin = 1;
#10 a = 24872; b = 2863; cin = 1;
#10 a = 61209; b = 56617; cin = 1;
#10 a = 11193; b = 40801; cin = 0;
#10 a = 56238; b = 50615; cin = 1;
#10 a = 47521; b = 14067; cin = 0;
#10 a = 13570; b = 47046; cin = 1;
#10 a = 68408; b = 34512; cin = 1;
#10 a = 30567; b = 29161; cin = 0;
#10 a = 43130; b = 53394; cin = 0;
#10 a = 15808; b = 60686; cin = 0;
#10 a = 1029; b = 61910; cin = 1;
#10 a = 51587; b = 29471; cin = 0;
#10 a = 18894; b = 40664; cin = 0;
#10 a = 58260; b = 3255; cin = 1;
#10 a = 63895; b = 50776; cin = 0;
#10 a = 45551; b = 40698; cin = 0;
#10 a = 43493; b = 15458; cin = 0;
#10 a = 21492; b = 46026; cin = 1;
#10 a = 68661; b = 19156; cin = 0;
#10 a = 7221; b = 34964; cin = 0;
#10 a = 36227; b = 12345; cin = 0;
#10 a = 44448; b = 63932; cin = 1;
#10 a = 39287; b = 59179; cin = 1;
#10 a = 51279; b = 23791; cin = 0;
#10 a = 20238; b = 64039; cin = 0;
#10 a = 3264; b = 39590; cin = 1;
#10 a = 33336; b = 59435; cin = 1;
#10 a = 4272; b = 10928; cin = 1;
#10 a = 50722; b = 55941; cin = 1;
#10 a = 10566; b = 63162; cin = 1;
#10 a = 7448; b = 29389; cin = 1;
#10 a = 42592; b = 50189; cin = 1;
#10 a = 37207; b = 19476; cin = 0;
#10 a = 48838; b = 47107; cin = 0;
#10 a = 63725; b = 43697; cin = 1;
#10 a = 35739; b = 46961; cin = 1;
#10 a = 48452; b = 10297; cin = 1;
#10 a = 52976; b = 60922; cin = 1;
#10 a = 33525; b = 41644; cin = 0;
#10 a = 9583; b = 28562; cin = 0;
#10 a = 20604; b = 12362; cin = 1;
#10 a = 20323; b = 54954; cin = 0;
#10 a = 60327; b = 22161; cin = 1;
#10 a = 65861; b = 47351; cin = 0;
#10 a = 25187; b = 17428; cin = 0;
#10 a = 48552; b = 53168; cin = 1;
#10 a = 41508; b = 7972; cin = 1;
#10 a = 251; b = 60948; cin = 1;
#10 a = 39922; b = 826; cin = 1;
#10 a = 65534; b = 10409; cin = 1;
#10 a = 60660; b = 7365; cin = 1;
#10 a = 15175; b = 4041; cin = 1;
#10 a = 19879; b = 40720; cin = 0;
#10 a = 66764; b = 36581; cin = 1;
#10 a = 20757; b = 38121; cin = 0;
#10 a = 64799; b = 16673; cin = 0;
#10 a = 39450; b = 34533; cin = 0;
#10 a = 47103; b = 34784; cin = 1;
#10 a = 69326; b = 4706; cin = 1;
#10 a = 15897; b = 46592; cin = 0;
#10 a = 61030; b = 37252; cin = 1;
#10 a = 48525; b = 52427; cin = 0;
#10 a = 67326; b = 48659; cin = 0;
#10 a = 14640; b = 45423; cin = 0;
#10 a = 32954; b = 42532; cin = 1;
#10 a = 45048; b = 37331; cin = 0;
#10 a = 16662; b = 53134; cin = 0;
#10 a = 66248; b = 30237; cin = 0;
#10 a = 36783; b = 5916; cin = 1;
#10 a = 30848; b = 68165; cin = 1;
#10 a = 58970; b = 35548; cin = 0;
#10 a = 810; b = 60425; cin = 1;
#10 a = 63042; b = 57752; cin = 0;
#10 a = 49643; b = 2392; cin = 0;
#10 a = 49177; b = 11698; cin = 0;
#10 a = 63184; b = 33098; cin = 0;
#10 a = 47512; b = 49760; cin = 0;
#10 a = 19078; b = 46009; cin = 1;
#10 a = 49077; b = 59144; cin = 1;
#10 a = 60134; b = 19993; cin = 1;
#10 a = 47783; b = 55315; cin = 1;
#10 a = 49037; b = 32477; cin = 0;
#10 a = 32719; b = 25520; cin = 0;
#10 a = 65059; b = 51515; cin = 1;
#10 a = 49175; b = 7044; cin = 1;
#10 a = 52176; b = 228; cin = 0;
#10 a = 22508; b = 24092; cin = 0;
#10 a = 45974; b = 43171; cin = 1;
#10 a = 52381; b = 22248; cin = 0;
#10 a = 64705; b = 58734; cin = 1;
#10 a = 51546; b = 12869; cin = 0;
#10 a = 27583; b = 61907; cin = 0;
#10 a = 40397; b = 24626; cin = 0;
#10 a = 40964; b = 19685; cin = 1;
#10 a = 20275; b = 45213; cin = 1;
#10 a = 57636; b = 27389; cin = 1;
#10 a = 58096; b = 49897; cin = 1;
#10 a = 14669; b = 2223; cin = 0;
#10 a = 17250; b = 30956; cin = 0;
#10 a = 55328; b = 25661; cin = 0;
#10 a = 43399; b = 7207; cin = 0;
#10 a = 39490; b = 11142; cin = 1;
#10 a = 21706; b = 27892; cin = 1;
#10 a = 52146; b = 68856; cin = 0;
#10 a = 17749; b = 65483; cin = 1;
#10 a = 60396; b = 29471; cin = 0;
#10 a = 9623; b = 63920; cin = 1;
#10 a = 6590; b = 8589; cin = 0;
#10 a = 23081; b = 25839; cin = 1;
#10 a = 61819; b = 11168; cin = 0;
#10 a = 19292; b = 30919; cin = 0;
#10 a = 35986; b = 46761; cin = 0;
#10 a = 44587; b = 44819; cin = 0;
#10 a = 7814; b = 26965; cin = 0;
#10 a = 13430; b = 44714; cin = 1;
#10 a = 64260; b = 11462; cin = 1;
#10 a = 2478; b = 21085; cin = 1;
#10 a = 36946; b = 27676; cin = 0;
#10 a = 49988; b = 50757; cin = 1;
#10 a = 23987; b = 18928; cin = 1;
#10 a = 23648; b = 38220; cin = 1;
#10 a = 53220; b = 50558; cin = 0;
#10 a = 47582; b = 25145; cin = 0;
#10 a = 46189; b = 9311; cin = 1;
#10 a = 20003; b = 22742; cin = 0;
#10 a = 35653; b = 17002; cin = 0;
#10 a = 10774; b = 65832; cin = 0;
#10 a = 26167; b = 32778; cin = 0;
#10 a = 50149; b = 59119; cin = 1;
#10 a = 29970; b = 13106; cin = 1;
#10 a = 43664; b = 13106; cin = 0;
#10 a = 18277; b = 66326; cin = 0;
#10 a = 16003; b = 20261; cin = 0;
#10 a = 12197; b = 42802; cin = 1;
#10 a = 11709; b = 62805; cin = 1;
#10 a = 32287; b = 4810; cin = 1;
#10 a = 17975; b = 61936; cin = 0;
#10 a = 1101; b = 18103; cin = 0;
#10 a = 11903; b = 44604; cin = 1;
#10 a = 26166; b = 4575; cin = 0;
#10 a = 13006; b = 48239; cin = 0;
#10 a = 60770; b = 42868; cin = 1;
#10 a = 19092; b = 58871; cin = 0;
#10 a = 2560; b = 47421; cin = 0;
#10 a = 41692; b = 35482; cin = 1;
#10 a = 9917; b = 67769; cin = 0;
#10 a = 65145; b = 62096; cin = 0;
#10 a = 22557; b = 63198; cin = 0;
#10 a = 12747; b = 51453; cin = 0;
#10 a = 62057; b = 7620; cin = 1;
#10 a = 54473; b = 20626; cin = 0;
#10 a = 36347; b = 57748; cin = 0;
#10 a = 14548; b = 6840; cin = 0;
#10 a = 36658; b = 55753; cin = 1;
#10 a = 7922; b = 27445; cin = 1;
#10 a = 18344; b = 13714; cin = 0;
#10 a = 9928; b = 55211; cin = 0;
#10 a = 63448; b = 7768; cin = 0;
#10 a = 65072; b = 20516; cin = 0;
#10 a = 17653; b = 58925; cin = 0;
#10 a = 21160; b = 19750; cin = 0;
#10 a = 2907; b = 56097; cin = 0;
#10 a = 3873; b = 646; cin = 0;
#10 a = 63711; b = 13656; cin = 1;
#10 a = 7322; b = 67931; cin = 0;
#10 a = 32767; b = 16275; cin = 1;
#10 a = 55981; b = 2555; cin = 0;
#10 a = 1292; b = 66003; cin = 1;
#10 a = 56152; b = 37428; cin = 1;
#10 a = 22466; b = 31433; cin = 0;
#10 a = 66400; b = 52593; cin = 0;
#10 a = 37312; b = 55500; cin = 1;
#10 a = 65972; b = 35726; cin = 1;
#10 a = 31473; b = 29437; cin = 0;
#10 a = 52726; b = 13112; cin = 1;
#10 a = 7777; b = 45879; cin = 0;
#10 a = 22894; b = 31861; cin = 1;
#10 a = 23222; b = 9505; cin = 0;
#10 a = 31319; b = 65657; cin = 0;
#10 a = 12636; b = 64476; cin = 1;
#10 a = 52878; b = 60876; cin = 1;
#10 a = 66518; b = 4541; cin = 1;
#10 a = 42608; b = 513; cin = 1;
#10 a = 65695; b = 31986; cin = 1;
#10 a = 56087; b = 61065; cin = 1;
#10 a = 20762; b = 45194; cin = 0;
#10 a = 48064; b = 68088; cin = 1;
#10 a = 7921; b = 21310; cin = 0;
#10 a = 33782; b = 28982; cin = 0;
#10 a = 3422; b = 17970; cin = 0;
#10 a = 4496; b = 849; cin = 0;
#10 a = 58163; b = 43719; cin = 1;
#10 a = 3682; b = 62679; cin = 1;
#10 a = 8576; b = 58375; cin = 1;
#10 a = 65611; b = 20814; cin = 0;
#10 a = 42110; b = 17929; cin = 0;
#10 a = 64488; b = 65993; cin = 0;
#10 a = 1432; b = 50267; cin = 1;
#10 a = 17880; b = 60401; cin = 1;
#10 a = 29986; b = 63823; cin = 1;
#10 a = 59272; b = 68319; cin = 0;
#10 a = 33083; b = 32834; cin = 0;
#10 a = 57786; b = 36517; cin = 1;
#10 a = 59355; b = 21445; cin = 0;
#10 a = 22911; b = 63408; cin = 1;
#10 a = 47531; b = 35518; cin = 0;
#10 a = 23698; b = 6358; cin = 1;
#10 a = 44304; b = 7790; cin = 0;
#10 a = 16221; b = 25671; cin = 1;
#10 a = 63472; b = 32009; cin = 1;
#10 a = 35046; b = 21282; cin = 0;
#10 a = 7468; b = 30717; cin = 1;
#10 a = 23610; b = 64855; cin = 0;
#10 a = 32432; b = 54211; cin = 1;
#10 a = 29628; b = 53474; cin = 1;
#10 a = 23991; b = 7357; cin = 1;
#10 a = 59931; b = 31055; cin = 1;
#10 a = 68217; b = 5360; cin = 0;
#10 a = 56769; b = 67933; cin = 1;
#10 a = 12075; b = 61406; cin = 0;
#10 a = 31204; b = 2804; cin = 0;
#10 a = 25004; b = 10272; cin = 1;
#10 a = 51639; b = 33883; cin = 1;
#10 a = 44791; b = 66315; cin = 0;
#10 a = 35740; b = 25943; cin = 0;
#10 a = 20097; b = 49935; cin = 1;
#10 a = 16324; b = 16218; cin = 1;
#10 a = 18910; b = 60787; cin = 1;
#10 a = 5638; b = 47557; cin = 0;
#10 a = 64389; b = 35984; cin = 0;
#10 a = 15149; b = 67188; cin = 0;
#10 a = 9896; b = 22192; cin = 1;
#10 a = 35359; b = 3832; cin = 0;
#10 a = 32030; b = 24975; cin = 1;
#10 a = 12912; b = 37068; cin = 0;
#10 a = 47268; b = 57165; cin = 1;
#10 a = 65334; b = 49842; cin = 0;
#10 a = 44455; b = 68752; cin = 1;
#10 a = 5288; b = 50742; cin = 0;
#10 a = 34054; b = 45131; cin = 0;
#10 a = 30579; b = 36632; cin = 0;
#10 a = 29907; b = 22880; cin = 1;
#10 a = 39508; b = 58240; cin = 1;
#10 a = 12992; b = 20270; cin = 0;
#10 a = 29143; b = 9535; cin = 0;
#10 a = 1238; b = 33155; cin = 0;
#10 a = 69619; b = 28489; cin = 0;
#10 a = 60571; b = 49296; cin = 0;
#10 a = 65959; b = 30936; cin = 0;
#10 a = 25255; b = 41343; cin = 1;
#10 a = 66888; b = 1922; cin = 1;
#10 a = 35708; b = 8181; cin = 0;
#10 a = 26721; b = 24042; cin = 0;
#10 a = 44270; b = 13386; cin = 0;
#10 a = 40443; b = 42530; cin = 1;
#10 a = 50035; b = 20120; cin = 1;
#10 a = 23145; b = 66091; cin = 0;
#10 a = 22449; b = 56663; cin = 1;
#10 a = 20505; b = 52622; cin = 1;
#10 a = 45655; b = 54229; cin = 0;
#10 a = 45936; b = 27469; cin = 0;
#10 a = 35554; b = 63178; cin = 0;
#10 a = 1700; b = 66251; cin = 0;
#10 a = 2438; b = 40522; cin = 0;
#10 a = 69798; b = 57317; cin = 0;
#10 a = 6694; b = 37352; cin = 0;
#10 a = 46745; b = 36850; cin = 0;
#10 a = 45285; b = 35651; cin = 1;
#10 a = 69474; b = 56157; cin = 1;
#10 a = 54600; b = 31812; cin = 0;
#10 a = 11068; b = 54101; cin = 0;
#10 a = 15811; b = 19655; cin = 0;
#10 a = 5087; b = 67707; cin = 1;
#10 a = 18405; b = 46497; cin = 1;
#10 a = 45109; b = 46295; cin = 0;
#10 a = 20696; b = 29341; cin = 1;
#10 a = 16402; b = 6086; cin = 1;
#10 a = 54552; b = 27724; cin = 0;
#10 a = 9365; b = 27198; cin = 1;
#10 a = 16800; b = 58150; cin = 0;
#10 a = 31169; b = 45571; cin = 1;
#10 a = 26655; b = 37734; cin = 0;
#10 a = 61671; b = 42821; cin = 1;
#10 a = 22938; b = 61226; cin = 0;
#10 a = 24728; b = 36335; cin = 1;
#10 a = 13834; b = 57031; cin = 1;
#10 a = 16645; b = 49786; cin = 1;
#10 a = 32658; b = 34338; cin = 1;
#10 a = 60675; b = 43704; cin = 0;
#10 a = 4848; b = 36856; cin = 0;
#10 a = 27186; b = 68025; cin = 1;
#10 a = 9977; b = 24680; cin = 1;
#10 a = 58775; b = 62703; cin = 0;
#10 a = 35280; b = 15642; cin = 0;
#10 a = 58282; b = 16722; cin = 0;
#10 a = 10284; b = 6908; cin = 1;
#10 a = 15275; b = 23554; cin = 1;
#10 a = 2704; b = 32564; cin = 0;
#10 a = 17858; b = 69591; cin = 0;
#10 a = 36562; b = 4440; cin = 0;
#10 a = 43416; b = 7978; cin = 0;
#10 a = 2194; b = 17956; cin = 0;
#10 a = 68705; b = 53083; cin = 0;
#10 a = 38038; b = 18364; cin = 0;
#10 a = 68596; b = 52998; cin = 0;
#10 a = 41842; b = 63282; cin = 0;
#10 a = 2120; b = 8557; cin = 0;
#10 a = 58535; b = 11262; cin = 1;
#10 a = 32937; b = 5472; cin = 0;
#10 a = 27395; b = 42034; cin = 0;
#10 a = 58710; b = 15450; cin = 1;
#10 a = 18050; b = 63996; cin = 1;
#10 a = 48422; b = 62702; cin = 0;
#10 a = 1498; b = 30740; cin = 0;
#10 a = 62920; b = 5688; cin = 1;
#10 a = 24712; b = 47531; cin = 1;
#10 a = 39765; b = 26003; cin = 1;
#10 a = 54723; b = 14538; cin = 1;
#10 a = 8598; b = 23828; cin = 1;
#10 a = 32065; b = 51223; cin = 1;
#10 a = 36323; b = 16285; cin = 1;
#10 a = 48560; b = 34335; cin = 0;
#10 a = 55105; b = 12758; cin = 0;
#10 a = 44734; b = 60608; cin = 0;
#10 a = 52726; b = 29881; cin = 0;
#10 a = 20069; b = 30945; cin = 1;
#10 a = 27047; b = 710; cin = 0;
#10 a = 42582; b = 31786; cin = 1;
#10 a = 69379; b = 40384; cin = 1;
#10 a = 54352; b = 48801; cin = 0;
#10 a = 35007; b = 15125; cin = 0;
#10 a = 7464; b = 63685; cin = 1;
#10 a = 20270; b = 48791; cin = 1;
#10 a = 25778; b = 69877; cin = 0;
#10 a = 62026; b = 28955; cin = 1;
#10 a = 33963; b = 49025; cin = 0;
#10 a = 29782; b = 6072; cin = 1;
#10 a = 51605; b = 48654; cin = 1;
#10 a = 17966; b = 24385; cin = 1;
#10 a = 8155; b = 8737; cin = 1;
#10 a = 25919; b = 20096; cin = 0;
#10 a = 59969; b = 3912; cin = 1;
#10 a = 34707; b = 24183; cin = 0;
#10 a = 22202; b = 49961; cin = 1;
#10 a = 46658; b = 41988; cin = 1;
#10 a = 7347; b = 52303; cin = 0;
#10 a = 68982; b = 12085; cin = 0;
#10 a = 61327; b = 63690; cin = 0;
#10 a = 38162; b = 58008; cin = 1;
#10 a = 55381; b = 66163; cin = 0;
#10 a = 51402; b = 68435; cin = 0;
#10 a = 62548; b = 34756; cin = 0;
#10 a = 43732; b = 69463; cin = 1;
#10 a = 50058; b = 21666; cin = 1;
#10 a = 9910; b = 44676; cin = 1;
#10 a = 45069; b = 28376; cin = 0;
#10 a = 59253; b = 27358; cin = 1;
#10 a = 55861; b = 65037; cin = 0;
#10 a = 7475; b = 33199; cin = 0;
#10 a = 6178; b = 64932; cin = 0;
#10 a = 13618; b = 46335; cin = 1;
#10 a = 41154; b = 15235; cin = 1;
#10 a = 48954; b = 35319; cin = 1;
#10 a = 34586; b = 15378; cin = 1;
#10 a = 46531; b = 1640; cin = 1;
#10 a = 6816; b = 46709; cin = 1;
#10 a = 19404; b = 35962; cin = 1;
#10 a = 44077; b = 68175; cin = 0;
#10 a = 15145; b = 52002; cin = 1;
#10 a = 67870; b = 58180; cin = 0;
#10 a = 69462; b = 1798; cin = 1;
#10 a = 23137; b = 19304; cin = 0;
#10 a = 57920; b = 68258; cin = 0;
#10 a = 68519; b = 9196; cin = 0;
#10 a = 30784; b = 32079; cin = 0;
#10 a = 14078; b = 38895; cin = 1;
#10 a = 25747; b = 34651; cin = 1;
#10 a = 41127; b = 55081; cin = 0;
#10 a = 51543; b = 226; cin = 0;
#10 a = 1511; b = 44448; cin = 0;
#10 a = 62763; b = 43910; cin = 0;
#10 a = 30350; b = 43399; cin = 0;
#10 a = 13172; b = 31320; cin = 0;
#10 a = 7666; b = 29839; cin = 1;
#10 a = 17538; b = 36976; cin = 0;
#10 a = 5402; b = 51054; cin = 0;
#10 a = 63623; b = 6801; cin = 1;
#10 a = 64158; b = 47928; cin = 0;
#10 a = 39220; b = 5824; cin = 1;
#10 a = 66284; b = 53687; cin = 1;
#10 a = 57880; b = 46450; cin = 0;
#10 a = 51274; b = 6800; cin = 1;
#10 a = 40324; b = 66324; cin = 1;
#10 a = 27633; b = 50343; cin = 1;
#10 a = 490; b = 67881; cin = 1;
#10 a = 29074; b = 49636; cin = 1;
#10 a = 49258; b = 43259; cin = 0;
#10 a = 57742; b = 13770; cin = 1;
#10 a = 27658; b = 52990; cin = 1;
#10 a = 67801; b = 25627; cin = 0;
#10 a = 12393; b = 13507; cin = 0;
#10 a = 47247; b = 64782; cin = 0;
#10 a = 9148; b = 11458; cin = 0;
#10 a = 48722; b = 39091; cin = 1;
#10 a = 839; b = 39581; cin = 1;
#10 a = 13580; b = 45008; cin = 1;
#10 a = 7375; b = 24266; cin = 0;
#10 a = 30675; b = 58360; cin = 0;
#10 a = 31904; b = 62371; cin = 1;
#10 a = 38957; b = 60172; cin = 0;
#10 a = 6049; b = 48917; cin = 1;
#10 a = 19591; b = 26164; cin = 1;
#10 a = 62637; b = 35313; cin = 0;
#10 a = 32008; b = 60387; cin = 1;
#10 a = 51721; b = 61226; cin = 1;
#10 a = 45668; b = 4806; cin = 1;
#10 a = 65603; b = 58533; cin = 1;
#10 a = 58798; b = 19208; cin = 0;
#10 a = 65762; b = 51113; cin = 1;
#10 a = 32069; b = 66422; cin = 1;
#10 a = 24003; b = 2472; cin = 1;
#10 a = 29445; b = 68415; cin = 1;
#10 a = 6020; b = 61053; cin = 0;
#10 a = 40406; b = 69413; cin = 1;
#10 a = 43884; b = 51134; cin = 1;
#10 a = 63295; b = 3155; cin = 1;
#10 a = 34066; b = 45110; cin = 0;
#10 a = 5455; b = 33908; cin = 1;
#10 a = 11557; b = 29671; cin = 0;
#10 a = 33678; b = 61740; cin = 0;
#10 a = 68676; b = 15744; cin = 0;
#10 a = 36239; b = 21541; cin = 0;
#10 a = 29966; b = 3913; cin = 1;
#10 a = 35359; b = 44320; cin = 0;
#10 a = 7490; b = 64556; cin = 0;
#10 a = 40848; b = 57851; cin = 1;
#10 a = 55363; b = 68269; cin = 0;
#10 a = 34764; b = 50076; cin = 0;
#10 a = 9725; b = 61634; cin = 1;
#10 a = 12151; b = 1664; cin = 0;
#10 a = 57351; b = 340; cin = 0;
#10 a = 35024; b = 12931; cin = 1;
#10 a = 57464; b = 42898; cin = 0;
#10 a = 957; b = 54609; cin = 0;
#10 a = 60215; b = 38451; cin = 0;
#10 a = 6959; b = 9299; cin = 1;
#10 a = 3211; b = 41015; cin = 0;
#10 a = 44573; b = 52131; cin = 1;
#10 a = 49843; b = 38208; cin = 1;
#10 a = 14785; b = 26711; cin = 1;
#10 a = 64171; b = 14062; cin = 0;
#10 a = 59301; b = 49086; cin = 1;
#10 a = 5972; b = 12902; cin = 1;
#10 a = 2908; b = 13859; cin = 0;
#10 a = 44165; b = 50426; cin = 0;
#10 a = 9977; b = 33738; cin = 1;
#10 a = 9993; b = 13301; cin = 0;
#10 a = 54629; b = 57874; cin = 1;
#10 a = 9342; b = 14069; cin = 1;
#10 a = 48393; b = 5206; cin = 0;
#10 a = 19109; b = 69377; cin = 1;
#10 a = 60165; b = 58678; cin = 1;
#10 a = 20504; b = 41002; cin = 0;
#10 a = 94; b = 43911; cin = 1;
#10 a = 10644; b = 64428; cin = 0;
#10 a = 13294; b = 4405; cin = 0;
#10 a = 47948; b = 60750; cin = 1;
#10 a = 53616; b = 21732; cin = 1;
#10 a = 17768; b = 7426; cin = 0;
#10 a = 66479; b = 55820; cin = 1;
#10 a = 25550; b = 4929; cin = 0;
#10 a = 45035; b = 41446; cin = 1;
#10 a = 19958; b = 38302; cin = 1;
#10 a = 7784; b = 38396; cin = 0;
#10 a = 9470; b = 49041; cin = 0;
#10 a = 14286; b = 38687; cin = 0;
#10 a = 52840; b = 62987; cin = 0;
#10 a = 11047; b = 22956; cin = 0;
#10 a = 3480; b = 17076; cin = 1;
#10 a = 56334; b = 13555; cin = 1;
#10 a = 68043; b = 39105; cin = 0;
#10 a = 55482; b = 60492; cin = 0;
#10 a = 31599; b = 56803; cin = 0;
#10 a = 25070; b = 64587; cin = 1;
#10 a = 62453; b = 4057; cin = 0;
#10 a = 24263; b = 64695; cin = 1;
#10 a = 60479; b = 23887; cin = 1;
#10 a = 40150; b = 11286; cin = 1;
#10 a = 41552; b = 61118; cin = 1;
#10 a = 50381; b = 47453; cin = 0;
#10 a = 45030; b = 45496; cin = 0;
#10 a = 20960; b = 7330; cin = 0;
#10 a = 14688; b = 15281; cin = 1;
#10 a = 367; b = 40352; cin = 1;
#10 a = 47146; b = 32805; cin = 0;
#10 a = 2966; b = 57068; cin = 0;
#10 a = 43825; b = 23900; cin = 1;
#10 a = 7672; b = 40402; cin = 0;
#10 a = 40827; b = 11954; cin = 0;
#10 a = 44706; b = 62336; cin = 1;
#10 a = 38493; b = 13718; cin = 0;
#10 a = 47737; b = 34679; cin = 0;
#10 a = 47473; b = 25719; cin = 0;
#10 a = 34013; b = 26086; cin = 0;
#10 a = 61492; b = 3232; cin = 1;
#10 a = 23028; b = 52550; cin = 1;
#10 a = 25612; b = 26376; cin = 1;
#10 a = 52084; b = 10400; cin = 1;
#10 a = 66194; b = 51228; cin = 0;
#10 a = 25070; b = 2286; cin = 0;
#10 a = 7752; b = 17131; cin = 0;
#10 a = 12282; b = 64868; cin = 1;
#10 a = 24142; b = 42342; cin = 1;
#10 a = 27636; b = 52707; cin = 1;
#10 a = 25130; b = 20551; cin = 0;
#10 a = 8133; b = 19931; cin = 0;
#10 a = 48205; b = 45544; cin = 0;
#10 a = 18528; b = 3980; cin = 1;
#10 a = 29254; b = 174; cin = 1;
#10 a = 51934; b = 1596; cin = 1;
#10 a = 43302; b = 9348; cin = 1;
#10 a = 48388; b = 67982; cin = 1;
#10 a = 64506; b = 22125; cin = 1;
#10 a = 59991; b = 26113; cin = 0;
#10 a = 34266; b = 51244; cin = 1;
#10 a = 11774; b = 35729; cin = 1;
#10 a = 18185; b = 13934; cin = 1;
#10 a = 27323; b = 8815; cin = 1;
#10 a = 510; b = 38069; cin = 1;
#10 a = 47629; b = 66355; cin = 1;
#10 a = 27035; b = 39657; cin = 0;
#10 a = 23572; b = 18045; cin = 0;
#10 a = 61329; b = 12551; cin = 1;
#10 a = 1429; b = 48894; cin = 1;
#10 a = 16939; b = 59513; cin = 1;
#10 a = 6649; b = 47639; cin = 0;
#10 a = 62642; b = 65824; cin = 1;
#10 a = 531; b = 23148; cin = 0;
#10 a = 36048; b = 10; cin = 1;
#10 a = 48091; b = 47640; cin = 0;
#10 a = 38082; b = 51027; cin = 1;
#10 a = 37422; b = 4599; cin = 0;
#10 a = 34745; b = 65928; cin = 0;
#10 a = 30544; b = 43709; cin = 0;
#10 a = 52457; b = 60649; cin = 1;
#10 a = 31966; b = 43650; cin = 1;
#10 a = 23557; b = 12644; cin = 1;
#10 a = 29082; b = 13175; cin = 1;
#10 a = 43422; b = 25575; cin = 0;
#10 a = 25831; b = 3666; cin = 0;
#10 a = 50947; b = 18100; cin = 1;
#10 a = 45720; b = 55523; cin = 0;
#10 a = 58538; b = 20268; cin = 0;
#10 a = 36612; b = 27164; cin = 0;
#10 a = 63581; b = 9622; cin = 1;
#10 a = 56414; b = 17940; cin = 1;
#10 a = 26887; b = 17849; cin = 1;
#10 a = 63185; b = 46931; cin = 0;
#10 a = 5334; b = 20353; cin = 1;
#10 a = 17494; b = 22536; cin = 1;
#10 a = 53646; b = 3483; cin = 1;
#10 a = 825; b = 49203; cin = 0;
#10 a = 68955; b = 14094; cin = 0;
#10 a = 39366; b = 50706; cin = 1;
#10 a = 29838; b = 20639; cin = 1;
#10 a = 10959; b = 53406; cin = 1;
#10 a = 35730; b = 10293; cin = 1;
#10 a = 3145; b = 49830; cin = 0;
#10 a = 30087; b = 55165; cin = 0;
#10 a = 12604; b = 2659; cin = 0;
#10 a = 68787; b = 56306; cin = 0;
#10 a = 49422; b = 33483; cin = 1;
#10 a = 15581; b = 32439; cin = 1;
#10 a = 48359; b = 48157; cin = 0;
#10 a = 38302; b = 7995; cin = 1;
#10 a = 14219; b = 18954; cin = 1;
#10 a = 54429; b = 31036; cin = 1;
#10 a = 42488; b = 10533; cin = 1;
#10 a = 7478; b = 40620; cin = 0;
#10 a = 39174; b = 29576; cin = 0;
#10 a = 23407; b = 4715; cin = 0;
#10 a = 11123; b = 54137; cin = 1;
#10 a = 24394; b = 46070; cin = 0;
#10 a = 5408; b = 782; cin = 1;
#10 a = 59832; b = 15436; cin = 0;
#10 a = 64895; b = 6008; cin = 0;
#10 a = 53365; b = 60437; cin = 0;
#10 a = 52128; b = 9277; cin = 1;
#10 a = 30721; b = 63107; cin = 1;
#10 a = 40832; b = 8634; cin = 1;
#10 a = 53602; b = 8393; cin = 0;
#10 a = 29030; b = 19516; cin = 0;
#10 a = 61589; b = 20262; cin = 0;
#10 a = 9292; b = 2022; cin = 0;
#10 a = 5151; b = 61854; cin = 1;
#10 a = 9006; b = 56750; cin = 1;
#10 a = 8166; b = 40115; cin = 0;
#10 a = 14715; b = 22243; cin = 1;
#10 a = 55444; b = 29316; cin = 0;
#10 a = 43146; b = 46500; cin = 0;
#10 a = 60423; b = 30102; cin = 1;
#10 a = 58768; b = 59132; cin = 1;
#10 a = 41250; b = 27074; cin = 0;
#10 a = 46154; b = 36366; cin = 0;
#10 a = 51841; b = 17869; cin = 1;
#10 a = 49316; b = 26875; cin = 1;
#10 a = 52799; b = 11394; cin = 0;
#10 a = 46719; b = 26109; cin = 1;
#10 a = 2620; b = 11553; cin = 1;
#10 a = 21628; b = 31051; cin = 0;
#10 a = 49271; b = 67827; cin = 0;
#10 a = 15306; b = 56595; cin = 1;
#10 a = 23562; b = 4197; cin = 1;
#10 a = 5728; b = 50351; cin = 1;
#10 a = 36268; b = 32192; cin = 0;
#10 a = 58663; b = 57860; cin = 0;
#10 a = 67808; b = 40659; cin = 0;
#10 a = 23420; b = 17378; cin = 1;
#10 a = 1275; b = 66350; cin = 0;
#10 a = 31151; b = 17979; cin = 0;
#10 a = 61175; b = 67250; cin = 1;
#10 a = 4005; b = 58908; cin = 0;
#10 a = 5968; b = 12470; cin = 1;
#10 a = 11357; b = 64550; cin = 0;
#10 a = 53112; b = 7171; cin = 1;
#10 a = 19089; b = 65834; cin = 1;
#10 a = 11941; b = 63643; cin = 1;
#10 a = 62539; b = 63415; cin = 1;
#10 a = 69246; b = 64691; cin = 0;
#10 a = 63858; b = 25842; cin = 1;
#10 a = 65874; b = 63369; cin = 1;
#10 a = 65717; b = 67374; cin = 1;
#10 a = 28507; b = 49695; cin = 0;
#10 a = 65494; b = 61052; cin = 0;
#10 a = 59185; b = 20517; cin = 1;
#10 a = 15068; b = 15958; cin = 0;
#10 a = 28811; b = 27899; cin = 1;
#10 a = 59566; b = 66790; cin = 0;
#10 a = 37700; b = 66036; cin = 1;
#10 a = 58536; b = 36246; cin = 1;
#10 a = 50999; b = 32121; cin = 0;
#10 a = 17064; b = 4190; cin = 1;
#10 a = 42037; b = 9050; cin = 0;
#10 a = 32185; b = 50896; cin = 0;
#10 a = 16884; b = 40081; cin = 1;
#10 a = 8753; b = 31501; cin = 1;
#10 a = 66457; b = 36665; cin = 0;
#10 a = 508; b = 26231; cin = 0;
#10 a = 21623; b = 40283; cin = 0;
#10 a = 13780; b = 28819; cin = 1;
#10 a = 8132; b = 9818; cin = 0;
#10 a = 65852; b = 3234; cin = 0;
#10 a = 27299; b = 21624; cin = 0;
#10 a = 14793; b = 53809; cin = 1;
#10 a = 63340; b = 693; cin = 0;
#10 a = 38755; b = 9447; cin = 0;
#10 a = 30129; b = 52256; cin = 1;
#10 a = 49401; b = 52765; cin = 0;
#10 a = 41816; b = 4388; cin = 0;
#10 a = 30266; b = 64520; cin = 1;
#10 a = 31315; b = 49004; cin = 0;
#10 a = 40837; b = 44857; cin = 0;
#10 a = 54550; b = 48508; cin = 0;
#10 a = 53664; b = 39654; cin = 0;
#10 a = 33675; b = 9346; cin = 1;
#10 a = 30120; b = 48101; cin = 0;
#10 a = 58066; b = 8230; cin = 1;
#10 a = 52677; b = 33984; cin = 0;
#10 a = 3519; b = 5800; cin = 0;
#10 a = 64645; b = 12418; cin = 0;
#10 a = 60943; b = 43734; cin = 1;
#10 a = 67059; b = 60923; cin = 0;
#10 a = 6409; b = 45473; cin = 0;
#10 a = 37384; b = 5490; cin = 0;
#10 a = 52168; b = 15517; cin = 0;
#10 a = 43997; b = 45637; cin = 0;
#10 a = 21626; b = 10055; cin = 0;
#10 a = 5159; b = 62732; cin = 0;
#10 a = 17809; b = 66252; cin = 0;
#10 a = 11199; b = 37249; cin = 1;
#10 a = 45461; b = 28192; cin = 1;
#10 a = 58728; b = 25251; cin = 0;
#10 a = 46852; b = 31661; cin = 0;
#10 a = 36189; b = 69045; cin = 0;
#10 a = 65179; b = 27565; cin = 1;
#10 a = 33516; b = 47914; cin = 1;
#10 a = 49954; b = 69540; cin = 0;
#10 a = 50974; b = 51051; cin = 1;
#10 a = 15979; b = 68860; cin = 1;
#10 a = 33135; b = 56411; cin = 0;
#10 a = 62710; b = 8225; cin = 1;
#10 a = 42371; b = 66953; cin = 0;
#10 a = 12956; b = 20158; cin = 1;
#10 a = 29014; b = 56347; cin = 0;
#10 a = 3266; b = 27878; cin = 1;
#10 a = 16683; b = 61394; cin = 0;
#10 a = 28442; b = 41348; cin = 0;
#10 a = 3905; b = 68675; cin = 0;
#10 a = 18452; b = 61006; cin = 0;
#10 a = 5603; b = 24141; cin = 0;
#10 a = 53651; b = 63204; cin = 1;
#10 a = 36244; b = 11927; cin = 0;
#10 a = 44089; b = 24883; cin = 0;
#10 a = 59946; b = 30249; cin = 1;
#10 a = 4849; b = 33515; cin = 0;
#10 a = 23668; b = 26551; cin = 0;
#10 a = 66754; b = 54993; cin = 1;
#10 a = 39381; b = 35250; cin = 0;
#10 a = 63059; b = 30054; cin = 0;
#10 a = 61949; b = 35657; cin = 1;
#10 a = 47251; b = 19309; cin = 1;
#10 a = 17130; b = 55553; cin = 1;
#10 a = 53963; b = 5994; cin = 0;
#10 a = 17305; b = 65941; cin = 0;
#10 a = 13347; b = 47142; cin = 1;
#10 a = 37267; b = 47162; cin = 0;
#10 a = 52581; b = 43917; cin = 0;
#10 a = 15596; b = 13298; cin = 0;
#10 a = 23638; b = 52709; cin = 1;
#10 a = 22686; b = 44658; cin = 0;
#10 a = 22228; b = 21910; cin = 1;
#10 a = 14973; b = 15392; cin = 1;
#10 a = 65998; b = 45707; cin = 1;
#10 a = 1907; b = 63013; cin = 0;
#10 a = 38065; b = 52712; cin = 0;
#10 a = 14090; b = 19979; cin = 1;
#10 a = 40315; b = 48912; cin = 0;
#10 a = 27885; b = 40861; cin = 0;
#10 a = 27057; b = 64499; cin = 1;
#10 a = 9932; b = 17186; cin = 1;
#10 a = 4817; b = 15766; cin = 1;
#10 a = 19010; b = 30739; cin = 0;
#10 a = 41461; b = 3090; cin = 1;
#10 a = 23555; b = 4997; cin = 0;
#10 a = 47941; b = 19414; cin = 0;
#10 a = 49470; b = 33504; cin = 1;
#10 a = 28161; b = 50171; cin = 0;
#10 a = 27121; b = 54408; cin = 1;
#10 a = 39379; b = 11466; cin = 0;
#10 a = 34346; b = 21398; cin = 0;
#10 a = 50323; b = 2567; cin = 0;
#10 a = 18211; b = 67930; cin = 0;
#10 a = 47843; b = 39391; cin = 0;
#10 a = 6830; b = 39298; cin = 1;
#10 a = 51535; b = 63592; cin = 1;
#10 a = 8951; b = 43062; cin = 1;
#10 a = 56347; b = 47575; cin = 1;
#10 a = 35359; b = 4696; cin = 1;
#10 a = 8880; b = 20427; cin = 1;
#10 a = 23252; b = 54773; cin = 0;
#10 a = 31163; b = 11448; cin = 1;
#10 a = 54839; b = 29659; cin = 1;
#10 a = 15607; b = 7502; cin = 1;
#10 a = 25817; b = 60685; cin = 1;
#10 a = 41024; b = 42220; cin = 1;
#10 a = 51997; b = 51171; cin = 1;
#10 a = 2827; b = 13870; cin = 0;
#10 a = 3828; b = 49229; cin = 0;
#10 a = 59237; b = 34461; cin = 1;
#10 a = 56113; b = 34066; cin = 0;
#10 a = 50739; b = 41581; cin = 1;
#10 a = 24284; b = 2772; cin = 0;
#10 a = 65760; b = 18380; cin = 1;
#10 a = 6627; b = 20549; cin = 0;
#10 a = 9496; b = 61574; cin = 0;
#10 a = 29606; b = 19923; cin = 1;
#10 a = 69129; b = 22750; cin = 0;
#10 a = 62580; b = 26578; cin = 1;
#10 a = 37078; b = 15816; cin = 1;
#10 a = 32004; b = 48281; cin = 1;
#10 a = 11702; b = 5372; cin = 0;
#10 a = 49201; b = 29656; cin = 0;
#10 a = 22712; b = 1768; cin = 0;
#10 a = 3725; b = 54747; cin = 0;
#10 a = 21775; b = 64244; cin = 0;
#10 a = 12045; b = 23850; cin = 1;
#10 a = 29838; b = 69331; cin = 0;
#10 a = 61502; b = 38263; cin = 0;
#10 a = 48748; b = 5342; cin = 0;
#10 a = 46807; b = 37346; cin = 1;
#10 a = 32580; b = 25400; cin = 1;
#10 a = 36286; b = 50954; cin = 0;
#10 a = 66412; b = 3666; cin = 0;
#10 a = 21271; b = 7391; cin = 0;
#10 a = 43031; b = 5518; cin = 0;
#10 a = 32717; b = 17563; cin = 0;
#10 a = 65974; b = 23753; cin = 1;
#10 a = 4686; b = 61608; cin = 1;
#10 a = 39977; b = 16708; cin = 1;
#10 a = 21083; b = 63515; cin = 1;
#10 a = 3175; b = 26095; cin = 1;
#10 a = 14286; b = 38733; cin = 1;
#10 a = 7758; b = 35145; cin = 1;
#10 a = 26647; b = 32768; cin = 0;
#10 a = 6635; b = 5799; cin = 0;
#10 a = 4515; b = 14868; cin = 1;
#10 a = 48949; b = 57195; cin = 1;
#10 a = 46362; b = 61881; cin = 1;
#10 a = 34743; b = 31858; cin = 1;
#10 a = 52114; b = 29294; cin = 0;
#10 a = 59535; b = 32469; cin = 1;
#10 a = 68709; b = 23107; cin = 0;
#10 a = 12484; b = 30866; cin = 1;
#10 a = 6278; b = 33865; cin = 0;
#10 a = 53814; b = 40500; cin = 1;
#10 a = 60517; b = 21367; cin = 0;
#10 a = 37486; b = 316; cin = 1;
#10 a = 38209; b = 23030; cin = 0;
#10 a = 30540; b = 57774; cin = 1;
#10 a = 15931; b = 16240; cin = 1;
#10 a = 64837; b = 52128; cin = 0;
#10 a = 46190; b = 50837; cin = 1;
#10 a = 66276; b = 39673; cin = 1;
#10 a = 51508; b = 22303; cin = 0;
#10 a = 45860; b = 6118; cin = 0;
#10 a = 22363; b = 42987; cin = 1;
#10 a = 13735; b = 10473; cin = 1;
	end
endmodule

module pfa(p, g, s, a, b, cin);
   output p, g, s;
   input a, b, cin;
   
   xor (s, a, b, cin);
   xor (p, a, b);
   and (g, a, b);
endmodule

//cla module 4 bit
module cla(p_up, g_up, cout, p, g, cin);
	output p_up, g_up;
	output[3:0] cout;
	input[3:0] p, g;
	input cin;
	
   //assign p_up = &(p);
   and  (p_up, p);
   wire p3g2, p3p2g1, p3p2p1g0, p3p2p1p0cin;
   
   and (p3g2,p[3],g[2]);
   and (p3p2g1,p[3],p[2],g[1]);
   and (p3p2p1g0,p[3],p[2],p[1],g[0]);
   
   and (p3p2p1p0cin,p[3],p[2],p[1],p[0],cin);
   
   //assign g_up = g[3] | p[3]&g[2] | p[3]&p[2]&g[1] | p[3]&p[2]&p[1]&g[0];
   or  (g_up,g[3],p3g2,p3p2g1,p3p2p1g0);
   
   //assign cout[3] = g[3] | p[3]&g[2] | p[3]&p[2]&g[1] | p[3]&p[2]&p[1]&g[0] | p[3]&p[2]&p[1]&p[0]&cin;
   or (cout[3],g[3],p3g2,p3p2g1,p3p2p1g0,p3p2p1p0cin);
   
   wire p2g1,p2p1g0,p2p1p0cin,p1g0,p1p0cin,p0cin;
   
   and (p2g1,p[2],g[1]);
   and (p2p1g0,p[2],p[1],g[0]);
   and (p2p1p0cin,p[2],p[1],p[0],cin);
   and (p1g0,p[1],g[0]);
   and (p1p0cin,p[1],p[0],cin);
   and (p0cin,p[0],cin);
   
   //assign cout[2] = g[2] | p[2]&g[1] | p[2]&p[1]&g[0] | p[2]&p[1]&p[0]&cin;
   or (cout[2], g[2],p2g1,p2p1g0,p2p1p0cin);
   
   //assign cout[1] = g[1] | p[1]&g[0] | p[1]&p[0]&cin;
   or (cout[1],g[1],p1g0,p1p0cin);
   
   //assign cout[0] = g[0] | p[0]&cin;
   or  (cout[0],g[0],p0cin);
endmodule

//put the cla and  adders together to make them easier to merge
module adder4_cla(cout, s, p_up, g_up, a, b, cin);
	output cout, p_up, g_up;
	output[3:0] s;
	input[3:0] a, b;
	input cin;

   wire [3:0] p,g;
   wire [3:0] carry;
   
   pfa add0(p[0], g[0], s[0], a[0], b[0], cin);
   pfa add1(p[1], g[1], s[1], a[1], b[1], carry[0]);
   pfa add2(p[2], g[2], s[2], a[2], b[2], carry[1]);
   pfa add3(p[3], g[3], s[3], a[3], b[3], carry[2]);

   cla localcla(p_up, g_up, carry, p, g, cin);
   assign cout = carry[3];
endmodule

module add16(cout, s, p_up, g_up, a, b, cin);
	output cout, p_up, g_up;
	output[15:0] s;
	input[15:0] a,b;
	input cin;
	wire [3:0] carry, p, g;
	
   adder4_cla add1 (carry[0], s[3:0], p[0], g[0], a[3:0], b[3:0], cin);
   adder4_cla add2 (carry[1], s[7:4], p[1], g[1], a[7:4], b[7:4], carry[0]);
   adder4_cla add3 (carry[2], s[11:8], p[2], g[2], a[11:8], b[11:8], carry[1]);
   adder4_cla add4 (cout, s[15:12], p[3], g[3], a[15:12], b[15:12], carry[2]);
endmodule
